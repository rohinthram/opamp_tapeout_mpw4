magic
tech sky130A
timestamp 1640402886
<< nwell >>
rect -52 244 1098 6720
<< nmos >>
rect 77 12 177 191
rect 507 10 607 189
rect -83 -2092 17 -1091
rect 278 -2232 378 -230
rect 1249 -2149 1349 4140
<< pmos >>
rect 77 306 177 1307
rect 506 306 606 1307
rect 862 304 962 6593
<< ndiff >>
rect -617 1596 -590 1603
rect -617 1579 -612 1596
rect -595 1579 -590 1596
rect -617 1572 -590 1579
rect -541 1582 -514 1589
rect -541 1565 -536 1582
rect -519 1565 -514 1582
rect -541 1558 -514 1565
rect -617 -927 -590 -920
rect -617 -944 -612 -927
rect -595 -944 -590 -927
rect -617 -951 -590 -944
rect -469 1585 -442 1592
rect -469 1568 -464 1585
rect -447 1568 -442 1585
rect -469 1561 -442 1568
rect -348 1576 -321 1583
rect -348 1559 -343 1576
rect -326 1559 -321 1576
rect -348 1552 -321 1559
rect -541 -941 -514 -934
rect -541 -958 -536 -941
rect -519 -958 -514 -941
rect -541 -965 -514 -958
rect -469 -938 -442 -931
rect -469 -955 -464 -938
rect -447 -955 -442 -938
rect -469 -962 -442 -955
rect 1143 3979 1249 4140
rect 1143 3915 1166 3979
rect 1228 3915 1249 3979
rect 1143 3857 1249 3915
rect 1144 3479 1249 3857
rect 1144 3415 1166 3479
rect 1228 3415 1249 3479
rect 1144 2979 1249 3415
rect 1144 2915 1166 2979
rect 1228 2915 1249 2979
rect 1144 2479 1249 2915
rect 1144 2415 1166 2479
rect 1228 2415 1249 2479
rect 1144 1979 1249 2415
rect 1144 1915 1166 1979
rect 1228 1915 1249 1979
rect 1144 1479 1249 1915
rect 1144 1415 1166 1479
rect 1228 1415 1249 1479
rect 1144 979 1249 1415
rect 1144 915 1166 979
rect 1228 915 1249 979
rect 1144 479 1249 915
rect 1144 415 1166 479
rect 1228 415 1249 479
rect -25 170 77 191
rect -25 122 -6 170
rect 38 122 77 170
rect -25 83 77 122
rect -25 35 -5 83
rect 39 35 77 83
rect -25 12 77 35
rect 177 169 287 191
rect 177 121 214 169
rect 258 121 287 169
rect 177 65 287 121
rect 177 19 205 65
rect 251 19 287 65
rect 177 12 287 19
rect 405 170 507 189
rect 405 122 426 170
rect 470 122 507 170
rect 405 76 507 122
rect 405 28 425 76
rect 469 28 507 76
rect 405 10 507 28
rect 607 176 717 189
rect 607 118 639 176
rect 693 118 717 176
rect 607 77 717 118
rect 607 30 642 77
rect 688 30 717 77
rect 607 10 717 30
rect 1144 -21 1249 415
rect 1144 -85 1166 -21
rect 1228 -85 1249 -21
rect 173 -344 278 -230
rect 173 -393 192 -344
rect 255 -393 278 -344
rect 173 -529 278 -393
rect -349 -948 -322 -942
rect -349 -973 -322 -970
rect 173 -593 192 -529
rect 255 -593 278 -529
rect 173 -729 278 -593
rect 173 -793 192 -729
rect 255 -793 278 -729
rect 173 -929 278 -793
rect 173 -993 192 -929
rect 255 -993 278 -929
rect -188 -1213 -83 -1091
rect -188 -1259 -158 -1213
rect -110 -1259 -83 -1213
rect -188 -1413 -83 -1259
rect -188 -1459 -158 -1413
rect -110 -1459 -83 -1413
rect -188 -1613 -83 -1459
rect -188 -1659 -158 -1613
rect -110 -1659 -83 -1613
rect -188 -1813 -83 -1659
rect -188 -1859 -158 -1813
rect -110 -1859 -83 -1813
rect -188 -2013 -83 -1859
rect -188 -2059 -158 -2013
rect -110 -2059 -83 -2013
rect -188 -2092 -83 -2059
rect 17 -1210 130 -1091
rect 17 -1256 55 -1210
rect 103 -1256 130 -1210
rect 17 -1410 130 -1256
rect 17 -1456 55 -1410
rect 103 -1456 130 -1410
rect 17 -1610 130 -1456
rect 17 -1656 55 -1610
rect 103 -1656 130 -1610
rect 17 -1810 130 -1656
rect 17 -1856 55 -1810
rect 103 -1856 130 -1810
rect 17 -2010 130 -1856
rect 17 -2056 55 -2010
rect 103 -2056 130 -2010
rect 17 -2092 130 -2056
rect 173 -1129 278 -993
rect 173 -1193 192 -1129
rect 255 -1193 278 -1129
rect 173 -1329 278 -1193
rect 173 -1393 192 -1329
rect 255 -1393 278 -1329
rect 173 -1529 278 -1393
rect 173 -1593 192 -1529
rect 255 -1593 278 -1529
rect 173 -1729 278 -1593
rect 173 -1793 192 -1729
rect 255 -1793 278 -1729
rect 173 -1929 278 -1793
rect 173 -1993 192 -1929
rect 255 -1993 278 -1929
rect 173 -2129 278 -1993
rect 173 -2193 192 -2129
rect 255 -2193 278 -2129
rect 173 -2232 278 -2193
rect 378 -329 491 -230
rect 378 -393 405 -329
rect 468 -393 491 -329
rect 378 -529 491 -393
rect 378 -593 405 -529
rect 468 -593 491 -529
rect 378 -729 491 -593
rect 378 -793 405 -729
rect 468 -793 491 -729
rect 378 -929 491 -793
rect 378 -993 405 -929
rect 468 -993 491 -929
rect 378 -1129 491 -993
rect 378 -1193 405 -1129
rect 468 -1193 491 -1129
rect 378 -1329 491 -1193
rect 378 -1393 405 -1329
rect 468 -1393 491 -1329
rect 378 -1529 491 -1393
rect 378 -1593 405 -1529
rect 468 -1593 491 -1529
rect 378 -1729 491 -1593
rect 378 -1793 405 -1729
rect 468 -1793 491 -1729
rect 378 -1929 491 -1793
rect 378 -1993 405 -1929
rect 468 -1993 491 -1929
rect 378 -2129 491 -1993
rect 378 -2193 405 -2129
rect 468 -2193 491 -2129
rect 1144 -521 1249 -85
rect 1144 -585 1166 -521
rect 1228 -585 1249 -521
rect 1144 -1021 1249 -585
rect 1144 -1085 1166 -1021
rect 1228 -1085 1249 -1021
rect 1144 -1521 1249 -1085
rect 1144 -1585 1166 -1521
rect 1228 -1585 1249 -1521
rect 1144 -2021 1249 -1585
rect 1144 -2085 1166 -2021
rect 1228 -2085 1249 -2021
rect 1144 -2149 1249 -2085
rect 1349 3979 1462 4140
rect 1349 3915 1374 3979
rect 1436 3915 1462 3979
rect 1349 3479 1462 3915
rect 1349 3415 1374 3479
rect 1436 3415 1462 3479
rect 1349 2979 1462 3415
rect 1349 2915 1374 2979
rect 1436 2915 1462 2979
rect 1349 2479 1462 2915
rect 1349 2415 1374 2479
rect 1436 2415 1462 2479
rect 1349 1979 1462 2415
rect 1349 1915 1374 1979
rect 1436 1915 1462 1979
rect 1349 1479 1462 1915
rect 1349 1415 1374 1479
rect 1436 1415 1462 1479
rect 1349 979 1462 1415
rect 1349 915 1374 979
rect 1436 915 1462 979
rect 1349 479 1462 915
rect 1349 415 1374 479
rect 1436 415 1462 479
rect 1349 -21 1462 415
rect 1349 -85 1374 -21
rect 1436 -85 1462 -21
rect 1349 -521 1462 -85
rect 1349 -585 1374 -521
rect 1436 -585 1462 -521
rect 1349 -1021 1462 -585
rect 1349 -1085 1374 -1021
rect 1436 -1085 1462 -1021
rect 1349 -1521 1462 -1085
rect 1349 -1585 1374 -1521
rect 1436 -1585 1462 -1521
rect 1349 -2021 1462 -1585
rect 1349 -2085 1374 -2021
rect 1436 -2085 1462 -2021
rect 1349 -2149 1462 -2085
rect 378 -2232 491 -2193
<< pdiff >>
rect 756 6422 862 6593
rect 756 6349 776 6422
rect 844 6349 862 6422
rect 756 6310 862 6349
rect 757 5922 862 6310
rect 757 5849 776 5922
rect 844 5849 862 5922
rect 757 5422 862 5849
rect 757 5349 776 5422
rect 844 5349 862 5422
rect 757 4922 862 5349
rect 757 4849 776 4922
rect 844 4849 862 4922
rect 757 4422 862 4849
rect 757 4349 776 4422
rect 844 4349 862 4422
rect 757 3922 862 4349
rect 757 3849 776 3922
rect 844 3849 862 3922
rect 757 3422 862 3849
rect 757 3349 776 3422
rect 844 3349 862 3422
rect 757 2922 862 3349
rect 757 2849 776 2922
rect 844 2849 862 2922
rect 757 2422 862 2849
rect 757 2349 776 2422
rect 844 2349 862 2422
rect 757 1922 862 2349
rect 757 1849 776 1922
rect 844 1849 862 1922
rect 757 1422 862 1849
rect 757 1349 776 1422
rect 844 1349 862 1422
rect -28 1222 77 1307
rect -28 1150 -7 1222
rect 60 1150 77 1222
rect -28 1022 77 1150
rect -28 950 -7 1022
rect 60 950 77 1022
rect -28 822 77 950
rect -28 750 -7 822
rect 60 750 77 822
rect -28 622 77 750
rect -28 550 -7 622
rect 60 550 77 622
rect -28 422 77 550
rect -28 350 -7 422
rect 60 350 77 422
rect -28 306 77 350
rect 177 1222 290 1307
rect 177 1149 205 1222
rect 273 1149 290 1222
rect 177 1022 290 1149
rect 177 949 205 1022
rect 273 949 290 1022
rect 177 822 290 949
rect 177 749 205 822
rect 273 749 290 822
rect 177 622 290 749
rect 177 549 205 622
rect 273 549 290 622
rect 177 422 290 549
rect 177 349 205 422
rect 273 349 290 422
rect 177 306 290 349
rect 401 1222 506 1307
rect 401 1149 419 1222
rect 487 1149 506 1222
rect 401 1022 506 1149
rect 401 949 419 1022
rect 487 949 506 1022
rect 401 822 506 949
rect 401 749 419 822
rect 487 749 506 822
rect 401 622 506 749
rect 401 549 419 622
rect 487 549 506 622
rect 401 422 506 549
rect 401 349 419 422
rect 487 349 506 422
rect 401 306 506 349
rect 606 1222 719 1307
rect 606 1149 627 1222
rect 695 1149 719 1222
rect 606 1022 719 1149
rect 606 949 627 1022
rect 695 949 719 1022
rect 606 822 719 949
rect 606 749 627 822
rect 695 749 719 822
rect 606 622 719 749
rect 606 549 627 622
rect 695 549 719 622
rect 606 422 719 549
rect 606 349 627 422
rect 695 349 719 422
rect 606 306 719 349
rect 757 922 862 1349
rect 757 849 776 922
rect 844 849 862 922
rect 757 422 862 849
rect 757 349 776 422
rect 844 349 862 422
rect 757 304 862 349
rect 962 6422 1075 6593
rect 962 6349 982 6422
rect 1050 6349 1075 6422
rect 962 5922 1075 6349
rect 962 5849 982 5922
rect 1050 5849 1075 5922
rect 962 5422 1075 5849
rect 962 5349 982 5422
rect 1050 5349 1075 5422
rect 962 4922 1075 5349
rect 962 4849 982 4922
rect 1050 4849 1075 4922
rect 962 4422 1075 4849
rect 962 4349 982 4422
rect 1050 4349 1075 4422
rect 962 3922 1075 4349
rect 962 3849 982 3922
rect 1050 3849 1075 3922
rect 962 3422 1075 3849
rect 962 3349 982 3422
rect 1050 3349 1075 3422
rect 962 2922 1075 3349
rect 962 2849 982 2922
rect 1050 2849 1075 2922
rect 962 2422 1075 2849
rect 962 2349 982 2422
rect 1050 2349 1075 2422
rect 962 1922 1075 2349
rect 962 1849 982 1922
rect 1050 1849 1075 1922
rect 962 1422 1075 1849
rect 962 1349 982 1422
rect 1050 1349 1075 1422
rect 962 922 1075 1349
rect 962 849 982 922
rect 1050 849 1075 922
rect 962 422 1075 849
rect 962 349 982 422
rect 1050 349 1075 422
rect 962 304 1075 349
<< ndiffc >>
rect -612 1579 -595 1596
rect -536 1565 -519 1582
rect -612 -944 -595 -927
rect -464 1568 -447 1585
rect -343 1559 -326 1576
rect -536 -958 -519 -941
rect -464 -955 -447 -938
rect 1166 3915 1228 3979
rect 1166 3415 1228 3479
rect 1166 2915 1228 2979
rect 1166 2415 1228 2479
rect 1166 1915 1228 1979
rect 1166 1415 1228 1479
rect 1166 915 1228 979
rect 1166 415 1228 479
rect -6 122 38 170
rect -5 35 39 83
rect 214 121 258 169
rect 205 19 251 65
rect 426 122 470 170
rect 425 28 469 76
rect 639 118 693 176
rect 642 30 688 77
rect 1166 -85 1228 -21
rect 192 -393 255 -344
rect -349 -970 -324 -948
rect 192 -593 255 -529
rect 192 -793 255 -729
rect 192 -993 255 -929
rect -158 -1259 -110 -1213
rect -158 -1459 -110 -1413
rect -158 -1659 -110 -1613
rect -158 -1859 -110 -1813
rect -158 -2059 -110 -2013
rect 55 -1256 103 -1210
rect 55 -1456 103 -1410
rect 55 -1656 103 -1610
rect 55 -1856 103 -1810
rect 55 -2056 103 -2010
rect 192 -1193 255 -1129
rect 192 -1393 255 -1329
rect 192 -1593 255 -1529
rect 192 -1793 255 -1729
rect 192 -1993 255 -1929
rect 192 -2193 255 -2129
rect 405 -393 468 -329
rect 405 -593 468 -529
rect 405 -793 468 -729
rect 405 -993 468 -929
rect 405 -1193 468 -1129
rect 405 -1393 468 -1329
rect 405 -1593 468 -1529
rect 405 -1793 468 -1729
rect 405 -1993 468 -1929
rect 405 -2193 468 -2129
rect 1166 -585 1228 -521
rect 1166 -1085 1228 -1021
rect 1166 -1585 1228 -1521
rect 1166 -2085 1228 -2021
rect 1374 3915 1436 3979
rect 1374 3415 1436 3479
rect 1374 2915 1436 2979
rect 1374 2415 1436 2479
rect 1374 1915 1436 1979
rect 1374 1415 1436 1479
rect 1374 915 1436 979
rect 1374 415 1436 479
rect 1374 -85 1436 -21
rect 1374 -585 1436 -521
rect 1374 -1085 1436 -1021
rect 1374 -1585 1436 -1521
rect 1374 -2085 1436 -2021
<< pdiffc >>
rect 776 6349 844 6422
rect 776 5849 844 5922
rect 776 5349 844 5422
rect 776 4849 844 4922
rect 776 4349 844 4422
rect 776 3849 844 3922
rect 776 3349 844 3422
rect 776 2849 844 2922
rect 776 2349 844 2422
rect 776 1849 844 1922
rect 776 1349 844 1422
rect -7 1150 60 1222
rect -7 950 60 1022
rect -7 750 60 822
rect -7 550 60 622
rect -7 350 60 422
rect 205 1149 273 1222
rect 205 949 273 1022
rect 205 749 273 822
rect 205 549 273 622
rect 205 349 273 422
rect 419 1149 487 1222
rect 419 949 487 1022
rect 419 749 487 822
rect 419 549 487 622
rect 419 349 487 422
rect 627 1149 695 1222
rect 627 949 695 1022
rect 627 749 695 822
rect 627 549 695 622
rect 627 349 695 422
rect 776 849 844 922
rect 776 349 844 422
rect 982 6349 1050 6422
rect 982 5849 1050 5922
rect 982 5349 1050 5422
rect 982 4849 1050 4922
rect 982 4349 1050 4422
rect 982 3849 1050 3922
rect 982 3349 1050 3422
rect 982 2849 1050 2922
rect 982 2349 1050 2422
rect 982 1849 1050 1922
rect 982 1349 1050 1422
rect 982 849 1050 922
rect 982 349 1050 422
<< psubdiff >>
rect -734 1574 -658 1605
rect -734 1524 -722 1574
rect -673 1524 -658 1574
rect -734 -1203 -658 1524
rect 1577 4148 1655 4168
rect -734 -1235 -656 -1203
rect -734 -1293 -727 -1235
rect -664 -1293 -656 -1235
rect -734 -1321 -656 -1293
rect -733 -2345 -656 -1321
rect 1577 4108 1590 4148
rect 1641 4108 1655 4148
rect 1577 3648 1655 4108
rect 1577 3608 1590 3648
rect 1641 3608 1655 3648
rect 1577 3148 1655 3608
rect 1577 3108 1590 3148
rect 1641 3108 1655 3148
rect 1577 2648 1655 3108
rect 1577 2608 1590 2648
rect 1641 2608 1655 2648
rect 1577 2148 1655 2608
rect 1577 2108 1590 2148
rect 1641 2108 1655 2148
rect 1577 1648 1655 2108
rect 1577 1608 1590 1648
rect 1641 1608 1655 1648
rect 1577 1148 1655 1608
rect 1577 1108 1590 1148
rect 1641 1108 1655 1148
rect 1577 648 1655 1108
rect 1577 608 1590 648
rect 1641 608 1655 648
rect 1577 148 1655 608
rect 1577 108 1590 148
rect 1641 108 1655 148
rect 1577 -352 1655 108
rect 1577 -392 1590 -352
rect 1641 -392 1655 -352
rect 1577 -852 1655 -392
rect 1577 -892 1590 -852
rect 1641 -892 1655 -852
rect 1577 -1352 1655 -892
rect 1577 -1392 1590 -1352
rect 1641 -1392 1655 -1352
rect 1577 -1852 1655 -1392
rect 1577 -1892 1590 -1852
rect 1641 -1892 1655 -1852
rect 1577 -2345 1655 -1892
rect -733 -2352 1655 -2345
rect -733 -2354 1590 -2352
rect -733 -2393 -718 -2354
rect -669 -2358 1590 -2354
rect -669 -2393 -414 -2358
rect -733 -2397 -414 -2393
rect -365 -2360 1590 -2358
rect -365 -2397 -92 -2360
rect -733 -2400 -92 -2397
rect -43 -2400 408 -2360
rect 457 -2400 908 -2360
rect 957 -2400 1408 -2360
rect 1457 -2392 1590 -2360
rect 1641 -2392 1655 -2352
rect 1457 -2400 1655 -2392
rect -733 -2409 1655 -2400
<< nsubdiff >>
rect 640 6695 707 6696
rect 638 6683 1072 6695
rect 638 6636 647 6683
rect 694 6680 1072 6683
rect 694 6638 1009 6680
rect 1057 6638 1072 6680
rect 694 6636 1072 6638
rect 638 6630 1072 6636
rect 640 6250 707 6630
rect 640 6209 656 6250
rect 693 6209 707 6250
rect 640 5750 707 6209
rect 640 5709 656 5750
rect 693 5709 707 5750
rect 640 5642 707 5709
rect 640 5250 708 5642
rect 640 5209 656 5250
rect 693 5209 708 5250
rect 640 5049 708 5209
rect 641 4750 708 5049
rect 641 4709 656 4750
rect 693 4709 708 4750
rect 641 4364 708 4709
rect 641 4250 705 4364
rect 641 4209 656 4250
rect 693 4209 705 4250
rect 641 3750 705 4209
rect 641 3709 656 3750
rect 693 3709 705 3750
rect 641 3250 705 3709
rect 641 3209 656 3250
rect 693 3209 705 3250
rect 641 2750 705 3209
rect 641 2709 656 2750
rect 693 2709 705 2750
rect 641 2250 705 2709
rect 641 2209 656 2250
rect 693 2209 705 2250
rect 641 1750 705 2209
rect 641 1709 656 1750
rect 693 1709 705 1750
rect 641 1569 705 1709
rect 642 1501 705 1569
rect 642 1468 653 1501
rect 686 1468 705 1501
rect 642 1456 705 1468
rect 15 1446 705 1456
rect 15 1445 219 1446
rect 15 1412 33 1445
rect 66 1413 219 1445
rect 252 1413 404 1446
rect 437 1413 563 1446
rect 596 1413 705 1446
rect 66 1412 705 1413
rect 15 1401 705 1412
<< psubdiffcont >>
rect -722 1524 -673 1574
rect -727 -1293 -664 -1235
rect 1590 4108 1641 4148
rect 1590 3608 1641 3648
rect 1590 3108 1641 3148
rect 1590 2608 1641 2648
rect 1590 2108 1641 2148
rect 1590 1608 1641 1648
rect 1590 1108 1641 1148
rect 1590 608 1641 648
rect 1590 108 1641 148
rect 1590 -392 1641 -352
rect 1590 -892 1641 -852
rect 1590 -1392 1641 -1352
rect 1590 -1892 1641 -1852
rect -718 -2393 -669 -2354
rect -414 -2397 -365 -2358
rect -92 -2400 -43 -2360
rect 408 -2400 457 -2360
rect 908 -2400 957 -2360
rect 1408 -2400 1457 -2360
rect 1590 -2392 1641 -2352
<< nsubdiffcont >>
rect 647 6636 694 6683
rect 1009 6638 1057 6680
rect 656 6209 693 6250
rect 656 5709 693 5750
rect 656 5209 693 5250
rect 656 4709 693 4750
rect 656 4209 693 4250
rect 656 3709 693 3750
rect 656 3209 693 3250
rect 656 2709 693 2750
rect 656 2209 693 2250
rect 656 1709 693 1750
rect 653 1468 686 1501
rect 33 1412 66 1445
rect 219 1413 252 1446
rect 404 1413 437 1446
rect 563 1413 596 1446
<< poly >>
rect 862 6593 962 6616
rect 77 1351 177 1364
rect 77 1345 115 1351
rect 75 1331 115 1345
rect 142 1345 177 1351
rect 142 1331 607 1345
rect 75 1316 607 1331
rect 77 1307 177 1316
rect 506 1307 606 1316
rect 77 260 177 306
rect 506 260 606 306
rect 1249 4140 1349 4163
rect 862 280 962 304
rect 862 257 887 280
rect 947 257 962 280
rect 862 245 962 257
rect 77 191 177 225
rect 507 189 607 223
rect 77 -13 177 12
rect 507 2 607 10
rect 77 -59 103 -13
rect 150 -59 177 -13
rect 77 -79 177 -59
rect 506 -52 607 2
rect 506 -87 535 -52
rect 575 -87 607 -52
rect 506 -110 607 -87
rect 278 -230 378 -205
rect -83 -1044 17 -1036
rect -83 -1072 -61 -1044
rect -2 -1072 17 -1044
rect -83 -1091 17 -1072
rect -83 -2270 17 -2092
rect 278 -2270 378 -2232
rect 1249 -2270 1349 -2149
rect -83 -2306 1349 -2270
<< polycont >>
rect 115 1331 142 1351
rect 887 257 947 280
rect 103 -59 150 -13
rect 535 -87 575 -52
rect -61 -1072 -2 -1044
<< ndiffres >>
rect -622 1603 -585 1605
rect -622 1572 -617 1603
rect -590 1572 -585 1603
rect -622 -564 -585 1572
rect -546 1589 -509 1606
rect -546 1558 -541 1589
rect -514 1558 -509 1589
rect -622 -920 -586 -564
rect -622 -951 -617 -920
rect -590 -951 -586 -920
rect -622 -957 -586 -951
rect -546 -578 -509 1558
rect -474 1592 -437 1609
rect -474 1561 -469 1592
rect -442 1561 -437 1592
rect -474 -575 -437 1561
rect -353 1583 -316 1587
rect -353 1552 -348 1583
rect -321 1552 -316 1583
rect -546 -934 -510 -578
rect -546 -965 -541 -934
rect -514 -965 -510 -934
rect -546 -971 -510 -965
rect -474 -931 -438 -575
rect -474 -962 -469 -931
rect -442 -962 -438 -931
rect -474 -968 -438 -962
rect -353 -584 -316 1552
rect -353 -942 -317 -584
rect -353 -973 -349 -942
rect -322 -948 -317 -942
rect -324 -970 -317 -948
rect -322 -973 -317 -970
rect -353 -979 -317 -973
<< locali >>
rect -28278 9959 -27733 9969
rect -54529 9659 -53982 9660
rect -54529 9029 -54516 9659
rect -53995 9029 -53982 9659
rect -28278 9366 -28266 9959
rect -27745 9366 -27733 9959
rect -28278 9356 -27733 9366
rect -2526 9453 -2057 9458
rect -54529 9028 -53982 9029
rect -2526 8968 -2516 9453
rect -2067 8968 -2057 9453
rect -2526 8963 -2057 8968
rect 25749 9451 26215 9462
rect 25749 8857 25757 9451
rect 26207 8857 26215 9451
rect 25749 8846 26215 8857
rect 46149 9416 46615 9427
rect 46149 8822 46157 9416
rect 46607 8822 46615 9416
rect 46149 8811 46615 8822
rect -54848 8292 -53656 8554
rect -54848 7662 -54479 8292
rect -53958 7662 -53656 8292
rect -54848 1850 -53656 7662
rect -28468 8180 -27546 8378
rect 704 8251 808 8252
rect -1638 8249 808 8251
rect -1881 8248 808 8249
rect -28468 7571 -28342 8180
rect -27654 7571 -27546 8180
rect -2700 8012 808 8248
rect -2700 7861 -2491 8012
rect -28468 3568 -27546 7571
rect -2699 7527 -2491 7861
rect -2042 7527 808 8012
rect -2699 7244 808 7527
rect -1881 7242 808 7244
rect 640 6695 707 6696
rect 725 6695 808 7242
rect 25501 8020 26467 8197
rect 25501 7426 25774 8020
rect 26224 7426 26467 8020
rect 638 6683 1072 6695
rect 638 6636 647 6683
rect 694 6680 1072 6683
rect 694 6638 1009 6680
rect 1057 6638 1072 6680
rect 694 6636 1072 6638
rect 638 6630 1072 6636
rect 640 6250 707 6630
rect 788 6433 833 6630
rect 767 6422 854 6433
rect 767 6349 776 6422
rect 844 6349 854 6422
rect 767 6341 854 6349
rect 973 6422 1060 6432
rect 973 6349 982 6422
rect 1050 6349 1060 6422
rect 973 6340 1060 6349
rect 640 6209 656 6250
rect 693 6209 707 6250
rect 640 5750 707 6209
rect 767 5922 854 5933
rect 767 5849 776 5922
rect 844 5849 854 5922
rect 767 5841 854 5849
rect 973 5922 1060 5932
rect 973 5849 982 5922
rect 1050 5849 1060 5922
rect 973 5840 1060 5849
rect 640 5709 656 5750
rect 693 5709 707 5750
rect 640 5642 707 5709
rect 640 5250 708 5642
rect 767 5422 854 5433
rect 767 5349 776 5422
rect 844 5349 854 5422
rect 767 5341 854 5349
rect 973 5422 1060 5432
rect 973 5349 982 5422
rect 1050 5349 1060 5422
rect 973 5340 1060 5349
rect 640 5209 656 5250
rect 693 5209 708 5250
rect 640 5049 708 5209
rect 641 4750 708 5049
rect 767 4922 854 4933
rect 767 4849 776 4922
rect 844 4849 854 4922
rect 767 4841 854 4849
rect 973 4922 1060 4932
rect 973 4849 982 4922
rect 1050 4849 1060 4922
rect 973 4840 1060 4849
rect 641 4709 656 4750
rect 693 4709 708 4750
rect 641 4364 708 4709
rect 767 4422 854 4433
rect 641 4250 705 4364
rect 767 4349 776 4422
rect 844 4349 854 4422
rect 767 4341 854 4349
rect 973 4428 1060 4432
rect 25501 4429 26467 7426
rect 25499 4428 26467 4429
rect 973 4422 26467 4428
rect 973 4349 982 4422
rect 1050 4349 26467 4422
rect 973 4344 26467 4349
rect 45901 7985 46864 8162
rect 45901 7391 46174 7985
rect 46624 7391 46864 7985
rect 45901 4792 46864 7391
rect 973 4340 1060 4344
rect 641 4209 656 4250
rect 693 4209 705 4250
rect 641 3750 705 4209
rect 1177 3993 1217 4344
rect 1577 4148 1655 4168
rect 1577 4108 1590 4148
rect 1641 4108 1655 4148
rect 1154 3979 1241 3993
rect 767 3922 854 3933
rect 767 3849 776 3922
rect 844 3849 854 3922
rect 767 3841 854 3849
rect 973 3922 1060 3932
rect 973 3849 982 3922
rect 1050 3849 1060 3922
rect 1154 3915 1166 3979
rect 1228 3915 1241 3979
rect 1154 3901 1241 3915
rect 1362 3979 1449 3993
rect 1362 3915 1374 3979
rect 1436 3915 1449 3979
rect 1362 3901 1449 3915
rect 973 3840 1060 3849
rect 641 3709 656 3750
rect 693 3709 705 3750
rect -28468 3431 -89 3568
rect -54849 1834 -53656 1850
rect -54849 1825 -195 1834
rect -54849 1796 -233 1825
rect -199 1796 -195 1825
rect -54849 1772 -195 1796
rect -54849 1743 -235 1772
rect -201 1743 -195 1772
rect -54849 1738 -195 1743
rect -54147 1734 -195 1738
rect -138 1776 -89 3431
rect -138 1744 -128 1776
rect -97 1744 -89 1776
rect -138 1734 -89 1744
rect 641 3250 705 3709
rect 1577 3648 1655 4108
rect 1577 3608 1590 3648
rect 1641 3608 1655 3648
rect 1154 3479 1241 3493
rect 767 3422 854 3433
rect 767 3349 776 3422
rect 844 3349 854 3422
rect 767 3341 854 3349
rect 973 3422 1060 3432
rect 973 3349 982 3422
rect 1050 3349 1060 3422
rect 1154 3415 1166 3479
rect 1228 3415 1241 3479
rect 1154 3401 1241 3415
rect 1362 3479 1449 3493
rect 1362 3415 1374 3479
rect 1436 3415 1449 3479
rect 1362 3401 1449 3415
rect 973 3340 1060 3349
rect 641 3209 656 3250
rect 693 3209 705 3250
rect 641 2750 705 3209
rect 1577 3148 1655 3608
rect 1577 3108 1590 3148
rect 1641 3108 1655 3148
rect 1154 2979 1241 2993
rect 767 2922 854 2933
rect 767 2849 776 2922
rect 844 2849 854 2922
rect 767 2841 854 2849
rect 973 2922 1060 2932
rect 973 2849 982 2922
rect 1050 2849 1060 2922
rect 1154 2915 1166 2979
rect 1228 2915 1241 2979
rect 1154 2901 1241 2915
rect 1362 2979 1449 2993
rect 1362 2915 1374 2979
rect 1436 2915 1449 2979
rect 1362 2901 1449 2915
rect 973 2840 1060 2849
rect 641 2709 656 2750
rect 693 2709 705 2750
rect 641 2250 705 2709
rect 1577 2648 1655 3108
rect 1577 2608 1590 2648
rect 1641 2608 1655 2648
rect 1154 2479 1241 2493
rect 767 2422 854 2433
rect 767 2349 776 2422
rect 844 2349 854 2422
rect 767 2341 854 2349
rect 973 2422 1060 2432
rect 973 2349 982 2422
rect 1050 2349 1060 2422
rect 1154 2415 1166 2479
rect 1228 2415 1241 2479
rect 1154 2401 1241 2415
rect 1362 2479 1449 2493
rect 1362 2415 1374 2479
rect 1436 2415 1449 2479
rect 1362 2401 1449 2415
rect 973 2340 1060 2349
rect 641 2209 656 2250
rect 693 2209 705 2250
rect 641 1750 705 2209
rect 1577 2148 1655 2608
rect 1577 2108 1590 2148
rect 1641 2108 1655 2148
rect 1154 1979 1241 1993
rect 767 1922 854 1933
rect 767 1849 776 1922
rect 844 1849 854 1922
rect 767 1841 854 1849
rect 973 1922 1060 1932
rect 973 1849 982 1922
rect 1050 1849 1060 1922
rect 1154 1915 1166 1979
rect 1228 1915 1241 1979
rect 1154 1901 1241 1915
rect 1362 1979 1449 1993
rect 1362 1915 1374 1979
rect 1436 1915 1449 1979
rect 1362 1901 1449 1915
rect 973 1840 1060 1849
rect 641 1709 656 1750
rect 693 1709 705 1750
rect -615 1645 56 1671
rect -615 1605 -593 1645
rect -472 1609 -438 1611
rect -544 1606 -510 1607
rect -734 1574 -658 1605
rect -734 1524 -722 1574
rect -673 1524 -658 1574
rect -620 1596 -585 1605
rect -620 1579 -612 1596
rect -595 1579 -585 1596
rect -620 1569 -585 1579
rect -619 1561 -585 1569
rect -544 1598 -509 1606
rect -472 1598 -437 1609
rect -544 1585 -437 1598
rect -544 1582 -464 1585
rect -544 1565 -536 1582
rect -519 1568 -464 1582
rect -447 1568 -437 1585
rect -353 1580 -316 1587
rect -519 1565 -437 1568
rect -544 1563 -437 1565
rect -544 1555 -509 1563
rect -472 1558 -437 1563
rect -543 1547 -509 1555
rect -471 1550 -437 1558
rect -405 1576 -316 1580
rect -405 1559 -343 1576
rect -326 1559 -316 1576
rect -405 1558 -316 1559
rect -734 -1203 -658 1524
rect -623 -927 -577 -906
rect -623 -944 -612 -927
rect -595 -938 -577 -927
rect -555 -938 -501 -920
rect -595 -941 -501 -938
rect -595 -944 -536 -941
rect -623 -958 -536 -944
rect -519 -958 -501 -941
rect -552 -977 -501 -958
rect -483 -938 -429 -917
rect -483 -955 -464 -938
rect -447 -955 -429 -938
rect -483 -966 -429 -955
rect -480 -978 -429 -966
rect -405 -978 -380 1558
rect -354 1550 -316 1558
rect 25 1456 56 1645
rect 641 1569 705 1709
rect 642 1501 705 1569
rect 642 1468 653 1501
rect 686 1468 705 1501
rect 1577 1648 1655 2108
rect 1577 1608 1590 1648
rect 1641 1608 1655 1648
rect 642 1456 705 1468
rect 15 1446 705 1456
rect 15 1445 219 1446
rect 15 1412 33 1445
rect 66 1413 219 1445
rect 252 1413 404 1446
rect 437 1413 563 1446
rect 596 1413 705 1446
rect 1154 1479 1241 1493
rect 66 1412 705 1413
rect 15 1401 705 1412
rect 767 1422 854 1433
rect 77 1351 177 1358
rect 77 1345 115 1351
rect -7 1331 115 1345
rect 142 1331 177 1351
rect -7 1315 177 1331
rect -7 1233 55 1315
rect 77 1314 177 1315
rect 209 1233 268 1401
rect 424 1233 482 1401
rect 767 1349 776 1422
rect 844 1349 854 1422
rect 767 1341 854 1349
rect 973 1422 1060 1432
rect 973 1349 982 1422
rect 1050 1349 1060 1422
rect 1154 1415 1166 1479
rect 1228 1415 1241 1479
rect 1154 1401 1241 1415
rect 1362 1479 1449 1493
rect 1362 1415 1374 1479
rect 1436 1415 1449 1479
rect 1362 1401 1449 1415
rect 973 1340 1060 1349
rect -16 1222 71 1233
rect -16 1150 -7 1222
rect 60 1150 71 1222
rect -16 1141 71 1150
rect 195 1222 282 1233
rect 195 1149 205 1222
rect 273 1149 282 1222
rect 195 1141 282 1149
rect 410 1222 497 1233
rect 410 1149 419 1222
rect 487 1149 497 1222
rect 410 1141 497 1149
rect 617 1222 704 1233
rect 617 1149 627 1222
rect 695 1149 704 1222
rect 617 1141 704 1149
rect 1577 1148 1655 1608
rect 1577 1108 1590 1148
rect 1641 1108 1655 1148
rect -16 1022 71 1033
rect -16 950 -7 1022
rect 60 950 71 1022
rect -16 941 71 950
rect 195 1022 282 1033
rect 195 949 205 1022
rect 273 949 282 1022
rect 195 941 282 949
rect 410 1022 497 1033
rect 410 949 419 1022
rect 487 949 497 1022
rect 410 941 497 949
rect 617 1022 704 1033
rect 617 949 627 1022
rect 695 949 704 1022
rect 617 941 704 949
rect 1154 979 1241 993
rect 767 922 854 933
rect 767 849 776 922
rect 844 849 854 922
rect 767 841 854 849
rect 973 922 1060 932
rect 973 849 982 922
rect 1050 849 1060 922
rect 1154 915 1166 979
rect 1228 915 1241 979
rect 1154 901 1241 915
rect 1362 979 1449 993
rect 1362 915 1374 979
rect 1436 915 1449 979
rect 1362 901 1449 915
rect 973 840 1060 849
rect -16 822 71 833
rect -16 750 -7 822
rect 60 750 71 822
rect -16 741 71 750
rect 195 822 282 833
rect 195 749 205 822
rect 273 749 282 822
rect 195 741 282 749
rect 410 822 497 833
rect 410 749 419 822
rect 487 749 497 822
rect 410 741 497 749
rect 617 822 704 833
rect 617 749 627 822
rect 695 749 704 822
rect 617 741 704 749
rect 1577 648 1655 1108
rect -16 622 71 633
rect -16 550 -7 622
rect 60 550 71 622
rect -16 541 71 550
rect 195 622 282 633
rect 195 549 205 622
rect 273 549 282 622
rect 195 541 282 549
rect 410 622 497 633
rect 410 549 419 622
rect 487 549 497 622
rect 410 541 497 549
rect 617 622 704 633
rect 617 549 627 622
rect 695 549 704 622
rect 617 541 704 549
rect 1577 608 1590 648
rect 1641 608 1655 648
rect 1154 479 1241 493
rect -16 422 71 433
rect -16 350 -7 422
rect 60 350 71 422
rect -16 341 71 350
rect 195 422 282 433
rect 195 349 205 422
rect 273 349 282 422
rect 195 341 282 349
rect 409 422 496 433
rect 409 349 419 422
rect 487 349 496 422
rect 409 341 496 349
rect 617 422 704 433
rect 617 349 627 422
rect 695 349 704 422
rect 617 341 704 349
rect 767 422 854 433
rect 767 349 776 422
rect 844 349 854 422
rect 767 341 854 349
rect 973 422 1060 432
rect 973 349 982 422
rect 1050 349 1060 422
rect 1154 415 1166 479
rect 1228 415 1241 479
rect 1154 401 1241 415
rect 1362 479 1449 493
rect 1362 415 1374 479
rect 1436 415 1449 479
rect 1362 401 1449 415
rect -6 180 40 341
rect 631 290 698 341
rect 973 340 1060 349
rect 862 290 962 299
rect 631 280 962 290
rect 631 257 887 280
rect 947 257 962 280
rect 631 256 962 257
rect -18 170 48 180
rect -18 122 -6 170
rect 38 122 48 170
rect -18 109 48 122
rect 202 169 268 180
rect 202 121 214 169
rect 258 121 268 169
rect 202 110 268 121
rect 412 170 478 178
rect 412 122 426 170
rect 470 122 478 170
rect 631 176 698 256
rect 862 245 962 256
rect 631 140 639 176
rect 412 107 478 122
rect 632 118 639 140
rect 693 118 698 176
rect 632 107 698 118
rect 1577 148 1655 608
rect 1577 108 1590 148
rect 1641 108 1655 148
rect -18 83 48 91
rect -18 35 -5 83
rect 39 35 48 83
rect -18 20 48 35
rect 190 76 266 80
rect 412 76 478 89
rect 190 65 425 76
rect 190 19 205 65
rect 251 28 425 65
rect 469 28 478 76
rect 251 19 478 28
rect 632 77 698 90
rect 632 30 642 77
rect 688 30 698 77
rect 632 19 698 30
rect 190 18 478 19
rect 190 16 472 18
rect 84 -13 169 1
rect 84 -59 103 -13
rect 150 -59 169 -13
rect 84 -78 169 -59
rect 190 -230 266 16
rect 1154 -21 1241 -7
rect 525 -52 585 -30
rect 525 -87 535 -52
rect 575 -87 585 -52
rect 525 -131 585 -87
rect 1154 -85 1166 -21
rect 1228 -85 1241 -21
rect 1154 -99 1241 -85
rect 1362 -21 1449 -7
rect 1362 -85 1374 -21
rect 1436 -85 1449 -21
rect 1362 -99 1449 -85
rect 525 -164 535 -131
rect 576 -164 585 -131
rect 525 -173 585 -164
rect 183 -344 265 -230
rect 183 -393 192 -344
rect 255 -393 265 -344
rect 183 -402 265 -393
rect 394 -329 476 -317
rect 394 -393 405 -329
rect 468 -393 476 -329
rect 394 -402 476 -393
rect 1577 -352 1655 108
rect 1577 -392 1590 -352
rect 1641 -392 1655 -352
rect 183 -529 265 -517
rect 183 -593 192 -529
rect 255 -593 265 -529
rect 183 -602 265 -593
rect 394 -529 476 -517
rect 394 -593 405 -529
rect 468 -593 476 -529
rect 394 -602 476 -593
rect 1154 -521 1241 -507
rect 1154 -585 1166 -521
rect 1228 -585 1241 -521
rect 1154 -599 1241 -585
rect 1362 -521 1449 -507
rect 1362 -585 1374 -521
rect 1436 -585 1449 -521
rect 1362 -599 1449 -585
rect 183 -729 265 -717
rect 183 -793 192 -729
rect 255 -793 265 -729
rect 183 -802 265 -793
rect 394 -729 476 -717
rect 394 -793 405 -729
rect 468 -793 476 -729
rect 394 -802 476 -793
rect 1577 -814 1655 -392
rect 45901 -814 46869 4792
rect 1577 -852 46869 -814
rect 1577 -892 1590 -852
rect 1641 -892 46869 -852
rect 183 -929 265 -917
rect -480 -998 -380 -978
rect -360 -948 -316 -943
rect -360 -970 -349 -948
rect -324 -970 -316 -948
rect -360 -979 -316 -970
rect -360 -1015 -110 -979
rect 183 -993 192 -929
rect 255 -993 265 -929
rect 183 -1002 265 -993
rect 394 -929 476 -917
rect 394 -993 405 -929
rect 468 -993 476 -929
rect 394 -1002 476 -993
rect -148 -1043 -110 -1015
rect 1154 -1021 1241 -1007
rect -83 -1043 17 -1040
rect -148 -1044 17 -1043
rect -148 -1072 -61 -1044
rect -2 -1072 17 -1044
rect -148 -1088 17 -1072
rect 1154 -1085 1166 -1021
rect 1228 -1085 1241 -1021
rect -148 -1201 -110 -1088
rect 1154 -1099 1241 -1085
rect 1362 -1021 1449 -1007
rect 1362 -1085 1374 -1021
rect 1436 -1085 1449 -1021
rect 1362 -1099 1449 -1085
rect 183 -1129 265 -1117
rect 183 -1193 192 -1129
rect 255 -1193 265 -1129
rect -734 -1235 -656 -1203
rect -734 -1293 -727 -1235
rect -664 -1293 -656 -1235
rect -171 -1213 -97 -1201
rect -171 -1259 -158 -1213
rect -110 -1259 -97 -1213
rect -171 -1273 -97 -1259
rect 42 -1210 116 -1197
rect 183 -1202 265 -1193
rect 394 -1129 476 -1117
rect 394 -1193 405 -1129
rect 468 -1193 476 -1129
rect 394 -1202 476 -1193
rect 1577 -1128 46869 -892
rect 42 -1256 55 -1210
rect 103 -1256 116 -1210
rect 42 -1270 116 -1256
rect -734 -1321 -656 -1293
rect -733 -2345 -656 -1321
rect 183 -1329 265 -1317
rect 183 -1393 192 -1329
rect 255 -1393 265 -1329
rect -171 -1413 -97 -1400
rect -171 -1459 -158 -1413
rect -110 -1459 -97 -1413
rect -171 -1473 -97 -1459
rect 42 -1410 116 -1397
rect 183 -1402 265 -1393
rect 394 -1329 476 -1317
rect 394 -1393 405 -1329
rect 468 -1393 476 -1329
rect 394 -1402 476 -1393
rect 1577 -1352 1655 -1128
rect 1577 -1392 1590 -1352
rect 1641 -1392 1655 -1352
rect 42 -1456 55 -1410
rect 103 -1456 116 -1410
rect 42 -1470 116 -1456
rect 183 -1529 265 -1517
rect 183 -1593 192 -1529
rect 255 -1593 265 -1529
rect -171 -1613 -97 -1600
rect -171 -1659 -158 -1613
rect -110 -1659 -97 -1613
rect -171 -1673 -97 -1659
rect 42 -1610 116 -1597
rect 183 -1602 265 -1593
rect 394 -1529 476 -1517
rect 394 -1593 405 -1529
rect 468 -1593 476 -1529
rect 394 -1602 476 -1593
rect 1154 -1521 1241 -1507
rect 1154 -1585 1166 -1521
rect 1228 -1585 1241 -1521
rect 1154 -1599 1241 -1585
rect 1362 -1521 1449 -1507
rect 1362 -1585 1374 -1521
rect 1436 -1585 1449 -1521
rect 1362 -1599 1449 -1585
rect 42 -1656 55 -1610
rect 103 -1656 116 -1610
rect 42 -1670 116 -1656
rect 183 -1729 265 -1717
rect 183 -1793 192 -1729
rect 255 -1793 265 -1729
rect -171 -1813 -97 -1800
rect -171 -1859 -158 -1813
rect -110 -1859 -97 -1813
rect -171 -1873 -97 -1859
rect 42 -1810 116 -1797
rect 183 -1802 265 -1793
rect 394 -1729 476 -1717
rect 394 -1793 405 -1729
rect 468 -1793 476 -1729
rect 394 -1802 476 -1793
rect 42 -1856 55 -1810
rect 103 -1856 116 -1810
rect 42 -1870 116 -1856
rect 1577 -1852 1655 -1392
rect 1577 -1892 1590 -1852
rect 1641 -1892 1655 -1852
rect 183 -1929 265 -1917
rect 183 -1993 192 -1929
rect 255 -1993 265 -1929
rect -173 -2013 -98 -2001
rect -173 -2059 -158 -2013
rect -110 -2059 -98 -2013
rect -173 -2075 -98 -2059
rect 40 -2010 115 -1998
rect 183 -2002 265 -1993
rect 394 -1929 476 -1917
rect 394 -1993 405 -1929
rect 468 -1993 476 -1929
rect 394 -2002 476 -1993
rect 40 -2056 55 -2010
rect 103 -2056 115 -2010
rect 40 -2072 115 -2056
rect 1154 -2021 1241 -2007
rect 49 -2345 111 -2072
rect 1154 -2085 1166 -2021
rect 1228 -2085 1241 -2021
rect 1154 -2099 1241 -2085
rect 1362 -2021 1449 -2007
rect 1362 -2085 1374 -2021
rect 1436 -2029 1449 -2021
rect 1577 -2029 1655 -1892
rect 1436 -2075 1655 -2029
rect 1436 -2085 1449 -2075
rect 1362 -2099 1449 -2085
rect 183 -2129 265 -2117
rect 183 -2193 192 -2129
rect 255 -2193 265 -2129
rect 183 -2202 265 -2193
rect 394 -2129 476 -2117
rect 394 -2193 405 -2129
rect 468 -2193 476 -2129
rect 394 -2202 476 -2193
rect 405 -2345 466 -2202
rect 1577 -2345 1655 -2075
rect -733 -2352 1655 -2345
rect -733 -2354 1590 -2352
rect -733 -2393 -718 -2354
rect -669 -2358 1590 -2354
rect -669 -2393 -414 -2358
rect -733 -2397 -414 -2393
rect -365 -2360 1590 -2358
rect -365 -2397 -92 -2360
rect -733 -2400 -92 -2397
rect -43 -2400 408 -2360
rect 457 -2400 908 -2360
rect 957 -2400 1408 -2360
rect 1457 -2392 1590 -2360
rect 1641 -2392 1655 -2352
rect 1457 -2400 1655 -2392
rect -733 -2409 1655 -2400
<< viali >>
rect -54516 9029 -53995 9659
rect -28266 9366 -27745 9959
rect -2516 8968 -2067 9453
rect 25757 8857 26207 9451
rect 46157 8822 46607 9416
rect -54479 7662 -53958 8292
rect -28342 7571 -27654 8180
rect -2491 7527 -2042 8012
rect 25774 7426 26224 8020
rect 46174 7391 46624 7985
rect -233 1796 -199 1825
rect -235 1743 -201 1772
rect -128 1744 -97 1776
rect 113 -50 136 -24
rect 535 -164 576 -131
<< metal1 >>
rect -54778 9659 -53685 10154
rect -54778 9645 -54516 9659
rect -53995 9645 -53685 9659
rect -54778 9043 -54525 9645
rect -53986 9043 -53685 9645
rect -54778 9029 -54516 9043
rect -53995 9029 -53685 9043
rect -54778 8292 -53685 9029
rect -54778 7662 -54479 8292
rect -53958 7662 -53685 8292
rect -54778 7256 -53685 7662
rect -28550 9964 -27507 10290
rect -28550 9361 -28275 9964
rect -27736 9361 -27507 9964
rect -28550 8180 -27507 9361
rect -28550 7571 -28342 8180
rect -27654 7571 -27507 8180
rect -2700 9453 -1770 10187
rect -2700 8968 -2516 9453
rect -2067 8968 -1770 9453
rect -2700 8012 -1770 8968
rect -2700 7861 -2491 8012
rect -28550 7398 -27507 7571
rect -2699 7527 -2491 7861
rect -2042 7527 -1770 8012
rect -2699 7288 -1770 7527
rect 25549 9455 26467 10051
rect 25549 9451 25761 9455
rect 26203 9451 26467 9455
rect 25549 8857 25757 9451
rect 26207 8857 26467 9451
rect 25549 8853 25761 8857
rect 26203 8853 26467 8857
rect 25549 8020 26467 8853
rect 25549 7426 25774 8020
rect 26224 7426 26467 8020
rect 25549 7166 26467 7426
rect 45949 9420 46864 10016
rect 45949 9416 46161 9420
rect 46603 9416 46864 9420
rect 45949 8822 46157 9416
rect 46607 8822 46864 9416
rect 45949 8818 46161 8822
rect 46603 8818 46864 8822
rect 45949 7985 46864 8818
rect 45949 7391 46174 7985
rect 46624 7391 46864 7985
rect 45949 7131 46864 7391
rect -244 1825 -195 1834
rect -244 1796 -233 1825
rect -199 1796 -195 1825
rect -244 1772 -195 1796
rect -244 1743 -235 1772
rect -201 1743 -195 1772
rect -244 -124 -195 1743
rect -138 1776 -89 1786
rect -138 1744 -128 1776
rect -97 1744 -89 1776
rect -138 -9 -89 1744
rect -138 -24 152 -9
rect -138 -50 113 -24
rect 136 -50 152 -24
rect -138 -60 152 -50
rect -244 -131 585 -124
rect -244 -164 535 -131
rect 576 -164 585 -131
rect -244 -173 585 -164
<< via1 >>
rect -54525 9043 -54516 9645
rect -54516 9043 -53995 9645
rect -53995 9043 -53986 9645
rect -28275 9959 -27736 9964
rect -28275 9366 -28266 9959
rect -28266 9366 -27745 9959
rect -27745 9366 -27736 9959
rect -28275 9361 -27736 9366
rect -2513 8973 -2070 9448
rect 25761 9451 26203 9455
rect 25761 8857 26203 9451
rect 25761 8853 26203 8857
rect 46161 9416 46603 9420
rect 46161 8822 46603 9416
rect 46161 8818 46603 8822
<< metal2 >>
rect -54778 9658 -53685 10154
rect -54778 9645 -54510 9658
rect -54001 9645 -53685 9658
rect -54778 9043 -54525 9645
rect -53986 9043 -53685 9645
rect -54778 9030 -54510 9043
rect -54001 9030 -53685 9043
rect -54778 7256 -53685 9030
rect -28550 9964 -27507 10290
rect -28550 9361 -28275 9964
rect -27736 9361 -27507 9964
rect -28550 7398 -27507 9361
rect -2700 9448 -1770 10187
rect -2700 9445 -2513 9448
rect -2070 9445 -1770 9448
rect -2700 8976 -2526 9445
rect -2057 8976 -1770 9445
rect -2700 8973 -2513 8976
rect -2070 8973 -1770 8976
rect -2700 7861 -1770 8973
rect -2699 7288 -1770 7861
rect 25549 9455 26467 10051
rect 25549 8853 25761 9455
rect 26203 8853 26467 9455
rect 25549 7166 26467 8853
rect 45949 9420 46864 10016
rect 45949 8818 46161 9420
rect 46603 8818 46864 9420
rect 45949 7131 46864 8818
<< via2 >>
rect -54510 9645 -54001 9658
rect -54510 9043 -54001 9645
rect -54510 9030 -54001 9043
rect -28260 9368 -27751 9957
rect -2526 8976 -2513 9445
rect -2513 8976 -2070 9445
rect -2070 8976 -2057 9445
rect 25768 8860 26196 9448
rect 46168 8825 46596 9413
<< metal3 >>
rect -54799 10917 -53659 11166
rect -54803 10791 -53659 10917
rect -54803 9658 -53662 10791
rect -28544 10692 -27473 11257
rect -2707 10837 -1737 11180
rect -28533 10290 -27477 10692
rect -54803 9189 -54510 9658
rect -54778 9030 -54510 9189
rect -54001 9189 -53662 9658
rect -28550 9957 -27477 10290
rect -28550 9368 -28260 9957
rect -27751 9816 -27477 9957
rect -27751 9368 -27507 9816
rect -54001 9030 -53685 9189
rect -54778 7256 -53685 9030
rect -28550 7398 -27507 9368
rect -2700 9667 -1739 10837
rect -2700 9445 -1770 9667
rect 24843 9516 26537 11079
rect 45765 10951 47464 11113
rect 45764 10930 47464 10951
rect -2700 8976 -2526 9445
rect -2057 8976 -1770 9445
rect 25516 9448 26467 9516
rect 25516 9212 25768 9448
rect -2700 7861 -1770 8976
rect -2699 7288 -1770 7861
rect 25549 8860 25768 9212
rect 26196 8860 26467 9448
rect 45764 9413 47458 10930
rect 45764 9388 46168 9413
rect 45916 9177 46168 9388
rect 25549 7166 26467 8860
rect 45949 8825 46168 9177
rect 46596 9388 47458 9413
rect 46596 8825 46864 9388
rect 45949 7131 46864 8825
<< labels >>
rlabel locali 835 6660 835 6660 1 vdd
rlabel locali 1192 4386 1192 4386 1 out
rlabel locali 705 -2384 705 -2384 1 vss
rlabel locali 551 -39 551 -39 1 in2
rlabel locali 124 -6 124 -6 1 in1
<< end >>
