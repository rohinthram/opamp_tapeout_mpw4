magic
tech sky130A
timestamp 1635438119
<< nwell >>
rect -54647 105229 -53497 111705
<< nmos >>
rect -54518 104997 -54418 105176
rect -54088 104995 -53988 105174
rect -54678 102893 -54578 103894
rect -54317 102753 -54217 104755
rect -53346 102836 -53246 109125
<< pmos >>
rect -54518 105291 -54418 106292
rect -54089 105291 -53989 106292
rect -53733 105289 -53633 111578
<< ndiff >>
rect -55212 106581 -55185 106588
rect -55212 106564 -55207 106581
rect -55190 106564 -55185 106581
rect -55212 106557 -55185 106564
rect -55136 106567 -55109 106574
rect -55136 106550 -55131 106567
rect -55114 106550 -55109 106567
rect -55136 106543 -55109 106550
rect -55212 104058 -55185 104065
rect -55212 104041 -55207 104058
rect -55190 104041 -55185 104058
rect -55212 104034 -55185 104041
rect -55064 106570 -55037 106577
rect -55064 106553 -55059 106570
rect -55042 106553 -55037 106570
rect -55064 106546 -55037 106553
rect -54943 106561 -54916 106568
rect -54943 106544 -54938 106561
rect -54921 106544 -54916 106561
rect -54943 106537 -54916 106544
rect -55136 104044 -55109 104051
rect -55136 104027 -55131 104044
rect -55114 104027 -55109 104044
rect -55136 104020 -55109 104027
rect -55064 104047 -55037 104054
rect -55064 104030 -55059 104047
rect -55042 104030 -55037 104047
rect -55064 104023 -55037 104030
rect -53452 108964 -53346 109125
rect -53452 108900 -53429 108964
rect -53367 108900 -53346 108964
rect -53452 108842 -53346 108900
rect -53451 108464 -53346 108842
rect -53451 108400 -53429 108464
rect -53367 108400 -53346 108464
rect -53451 107964 -53346 108400
rect -53451 107900 -53429 107964
rect -53367 107900 -53346 107964
rect -53451 107464 -53346 107900
rect -53451 107400 -53429 107464
rect -53367 107400 -53346 107464
rect -53451 106964 -53346 107400
rect -53451 106900 -53429 106964
rect -53367 106900 -53346 106964
rect -53451 106464 -53346 106900
rect -53451 106400 -53429 106464
rect -53367 106400 -53346 106464
rect -53451 105964 -53346 106400
rect -53451 105900 -53429 105964
rect -53367 105900 -53346 105964
rect -53451 105464 -53346 105900
rect -53451 105400 -53429 105464
rect -53367 105400 -53346 105464
rect -54620 105155 -54518 105176
rect -54620 105107 -54601 105155
rect -54557 105107 -54518 105155
rect -54620 105068 -54518 105107
rect -54620 105020 -54600 105068
rect -54556 105020 -54518 105068
rect -54620 104997 -54518 105020
rect -54418 105154 -54308 105176
rect -54418 105106 -54381 105154
rect -54337 105106 -54308 105154
rect -54418 105050 -54308 105106
rect -54418 105004 -54390 105050
rect -54344 105004 -54308 105050
rect -54418 104997 -54308 105004
rect -54190 105155 -54088 105174
rect -54190 105107 -54169 105155
rect -54125 105107 -54088 105155
rect -54190 105061 -54088 105107
rect -54190 105013 -54170 105061
rect -54126 105013 -54088 105061
rect -54190 104995 -54088 105013
rect -53988 105161 -53878 105174
rect -53988 105103 -53956 105161
rect -53902 105103 -53878 105161
rect -53988 105062 -53878 105103
rect -53988 105015 -53953 105062
rect -53907 105015 -53878 105062
rect -53988 104995 -53878 105015
rect -53451 104964 -53346 105400
rect -53451 104900 -53429 104964
rect -53367 104900 -53346 104964
rect -54422 104641 -54317 104755
rect -54422 104592 -54403 104641
rect -54340 104592 -54317 104641
rect -54422 104456 -54317 104592
rect -54944 104037 -54917 104043
rect -54944 104012 -54917 104015
rect -54422 104392 -54403 104456
rect -54340 104392 -54317 104456
rect -54422 104256 -54317 104392
rect -54422 104192 -54403 104256
rect -54340 104192 -54317 104256
rect -54422 104056 -54317 104192
rect -54422 103992 -54403 104056
rect -54340 103992 -54317 104056
rect -54783 103772 -54678 103894
rect -54783 103726 -54753 103772
rect -54705 103726 -54678 103772
rect -54783 103572 -54678 103726
rect -54783 103526 -54753 103572
rect -54705 103526 -54678 103572
rect -54783 103372 -54678 103526
rect -54783 103326 -54753 103372
rect -54705 103326 -54678 103372
rect -54783 103172 -54678 103326
rect -54783 103126 -54753 103172
rect -54705 103126 -54678 103172
rect -54783 102972 -54678 103126
rect -54783 102926 -54753 102972
rect -54705 102926 -54678 102972
rect -54783 102893 -54678 102926
rect -54578 103775 -54465 103894
rect -54578 103729 -54540 103775
rect -54492 103729 -54465 103775
rect -54578 103575 -54465 103729
rect -54578 103529 -54540 103575
rect -54492 103529 -54465 103575
rect -54578 103375 -54465 103529
rect -54578 103329 -54540 103375
rect -54492 103329 -54465 103375
rect -54578 103175 -54465 103329
rect -54578 103129 -54540 103175
rect -54492 103129 -54465 103175
rect -54578 102975 -54465 103129
rect -54578 102929 -54540 102975
rect -54492 102929 -54465 102975
rect -54578 102893 -54465 102929
rect -54422 103856 -54317 103992
rect -54422 103792 -54403 103856
rect -54340 103792 -54317 103856
rect -54422 103656 -54317 103792
rect -54422 103592 -54403 103656
rect -54340 103592 -54317 103656
rect -54422 103456 -54317 103592
rect -54422 103392 -54403 103456
rect -54340 103392 -54317 103456
rect -54422 103256 -54317 103392
rect -54422 103192 -54403 103256
rect -54340 103192 -54317 103256
rect -54422 103056 -54317 103192
rect -54422 102992 -54403 103056
rect -54340 102992 -54317 103056
rect -54422 102856 -54317 102992
rect -54422 102792 -54403 102856
rect -54340 102792 -54317 102856
rect -54422 102753 -54317 102792
rect -54217 104656 -54104 104755
rect -54217 104592 -54190 104656
rect -54127 104592 -54104 104656
rect -54217 104456 -54104 104592
rect -54217 104392 -54190 104456
rect -54127 104392 -54104 104456
rect -54217 104256 -54104 104392
rect -54217 104192 -54190 104256
rect -54127 104192 -54104 104256
rect -54217 104056 -54104 104192
rect -54217 103992 -54190 104056
rect -54127 103992 -54104 104056
rect -54217 103856 -54104 103992
rect -54217 103792 -54190 103856
rect -54127 103792 -54104 103856
rect -54217 103656 -54104 103792
rect -54217 103592 -54190 103656
rect -54127 103592 -54104 103656
rect -54217 103456 -54104 103592
rect -54217 103392 -54190 103456
rect -54127 103392 -54104 103456
rect -54217 103256 -54104 103392
rect -54217 103192 -54190 103256
rect -54127 103192 -54104 103256
rect -54217 103056 -54104 103192
rect -54217 102992 -54190 103056
rect -54127 102992 -54104 103056
rect -54217 102856 -54104 102992
rect -54217 102792 -54190 102856
rect -54127 102792 -54104 102856
rect -53451 104464 -53346 104900
rect -53451 104400 -53429 104464
rect -53367 104400 -53346 104464
rect -53451 103964 -53346 104400
rect -53451 103900 -53429 103964
rect -53367 103900 -53346 103964
rect -53451 103464 -53346 103900
rect -53451 103400 -53429 103464
rect -53367 103400 -53346 103464
rect -53451 102964 -53346 103400
rect -53451 102900 -53429 102964
rect -53367 102900 -53346 102964
rect -53451 102836 -53346 102900
rect -53246 108964 -53133 109125
rect -53246 108900 -53221 108964
rect -53159 108900 -53133 108964
rect -53246 108464 -53133 108900
rect -53246 108400 -53221 108464
rect -53159 108400 -53133 108464
rect -53246 107964 -53133 108400
rect -53246 107900 -53221 107964
rect -53159 107900 -53133 107964
rect -53246 107464 -53133 107900
rect -53246 107400 -53221 107464
rect -53159 107400 -53133 107464
rect -53246 106964 -53133 107400
rect -53246 106900 -53221 106964
rect -53159 106900 -53133 106964
rect -53246 106464 -53133 106900
rect -53246 106400 -53221 106464
rect -53159 106400 -53133 106464
rect -53246 105964 -53133 106400
rect -53246 105900 -53221 105964
rect -53159 105900 -53133 105964
rect -53246 105464 -53133 105900
rect -53246 105400 -53221 105464
rect -53159 105400 -53133 105464
rect -53246 104964 -53133 105400
rect -53246 104900 -53221 104964
rect -53159 104900 -53133 104964
rect -53246 104464 -53133 104900
rect -53246 104400 -53221 104464
rect -53159 104400 -53133 104464
rect -53246 103964 -53133 104400
rect -53246 103900 -53221 103964
rect -53159 103900 -53133 103964
rect -53246 103464 -53133 103900
rect -53246 103400 -53221 103464
rect -53159 103400 -53133 103464
rect -53246 102964 -53133 103400
rect -53246 102900 -53221 102964
rect -53159 102900 -53133 102964
rect -53246 102836 -53133 102900
rect -54217 102753 -54104 102792
<< pdiff >>
rect -53839 111407 -53733 111578
rect -53839 111334 -53819 111407
rect -53751 111334 -53733 111407
rect -53839 111295 -53733 111334
rect -53838 110907 -53733 111295
rect -53838 110834 -53819 110907
rect -53751 110834 -53733 110907
rect -53838 110407 -53733 110834
rect -53838 110334 -53819 110407
rect -53751 110334 -53733 110407
rect -53838 109907 -53733 110334
rect -53838 109834 -53819 109907
rect -53751 109834 -53733 109907
rect -53838 109407 -53733 109834
rect -53838 109334 -53819 109407
rect -53751 109334 -53733 109407
rect -53838 108907 -53733 109334
rect -53838 108834 -53819 108907
rect -53751 108834 -53733 108907
rect -53838 108407 -53733 108834
rect -53838 108334 -53819 108407
rect -53751 108334 -53733 108407
rect -53838 107907 -53733 108334
rect -53838 107834 -53819 107907
rect -53751 107834 -53733 107907
rect -53838 107407 -53733 107834
rect -53838 107334 -53819 107407
rect -53751 107334 -53733 107407
rect -53838 106907 -53733 107334
rect -53838 106834 -53819 106907
rect -53751 106834 -53733 106907
rect -53838 106407 -53733 106834
rect -53838 106334 -53819 106407
rect -53751 106334 -53733 106407
rect -54623 106207 -54518 106292
rect -54623 106135 -54602 106207
rect -54535 106135 -54518 106207
rect -54623 106007 -54518 106135
rect -54623 105935 -54602 106007
rect -54535 105935 -54518 106007
rect -54623 105807 -54518 105935
rect -54623 105735 -54602 105807
rect -54535 105735 -54518 105807
rect -54623 105607 -54518 105735
rect -54623 105535 -54602 105607
rect -54535 105535 -54518 105607
rect -54623 105407 -54518 105535
rect -54623 105335 -54602 105407
rect -54535 105335 -54518 105407
rect -54623 105291 -54518 105335
rect -54418 106207 -54305 106292
rect -54418 106134 -54390 106207
rect -54322 106134 -54305 106207
rect -54418 106007 -54305 106134
rect -54418 105934 -54390 106007
rect -54322 105934 -54305 106007
rect -54418 105807 -54305 105934
rect -54418 105734 -54390 105807
rect -54322 105734 -54305 105807
rect -54418 105607 -54305 105734
rect -54418 105534 -54390 105607
rect -54322 105534 -54305 105607
rect -54418 105407 -54305 105534
rect -54418 105334 -54390 105407
rect -54322 105334 -54305 105407
rect -54418 105291 -54305 105334
rect -54194 106207 -54089 106292
rect -54194 106134 -54176 106207
rect -54108 106134 -54089 106207
rect -54194 106007 -54089 106134
rect -54194 105934 -54176 106007
rect -54108 105934 -54089 106007
rect -54194 105807 -54089 105934
rect -54194 105734 -54176 105807
rect -54108 105734 -54089 105807
rect -54194 105607 -54089 105734
rect -54194 105534 -54176 105607
rect -54108 105534 -54089 105607
rect -54194 105407 -54089 105534
rect -54194 105334 -54176 105407
rect -54108 105334 -54089 105407
rect -54194 105291 -54089 105334
rect -53989 106207 -53876 106292
rect -53989 106134 -53968 106207
rect -53900 106134 -53876 106207
rect -53989 106007 -53876 106134
rect -53989 105934 -53968 106007
rect -53900 105934 -53876 106007
rect -53989 105807 -53876 105934
rect -53989 105734 -53968 105807
rect -53900 105734 -53876 105807
rect -53989 105607 -53876 105734
rect -53989 105534 -53968 105607
rect -53900 105534 -53876 105607
rect -53989 105407 -53876 105534
rect -53989 105334 -53968 105407
rect -53900 105334 -53876 105407
rect -53989 105291 -53876 105334
rect -53838 105907 -53733 106334
rect -53838 105834 -53819 105907
rect -53751 105834 -53733 105907
rect -53838 105407 -53733 105834
rect -53838 105334 -53819 105407
rect -53751 105334 -53733 105407
rect -53838 105289 -53733 105334
rect -53633 111407 -53520 111578
rect -53633 111334 -53613 111407
rect -53545 111334 -53520 111407
rect -53633 110907 -53520 111334
rect -53633 110834 -53613 110907
rect -53545 110834 -53520 110907
rect -53633 110407 -53520 110834
rect -53633 110334 -53613 110407
rect -53545 110334 -53520 110407
rect -53633 109907 -53520 110334
rect -53633 109834 -53613 109907
rect -53545 109834 -53520 109907
rect -53633 109407 -53520 109834
rect -53633 109334 -53613 109407
rect -53545 109334 -53520 109407
rect -53633 108907 -53520 109334
rect -53633 108834 -53613 108907
rect -53545 108834 -53520 108907
rect -53633 108407 -53520 108834
rect -53633 108334 -53613 108407
rect -53545 108334 -53520 108407
rect -53633 107907 -53520 108334
rect -53633 107834 -53613 107907
rect -53545 107834 -53520 107907
rect -53633 107407 -53520 107834
rect -53633 107334 -53613 107407
rect -53545 107334 -53520 107407
rect -53633 106907 -53520 107334
rect -53633 106834 -53613 106907
rect -53545 106834 -53520 106907
rect -53633 106407 -53520 106834
rect -53633 106334 -53613 106407
rect -53545 106334 -53520 106407
rect -53633 105907 -53520 106334
rect -53633 105834 -53613 105907
rect -53545 105834 -53520 105907
rect -53633 105407 -53520 105834
rect -53633 105334 -53613 105407
rect -53545 105334 -53520 105407
rect -53633 105289 -53520 105334
<< ndiffc >>
rect -55207 106564 -55190 106581
rect -55131 106550 -55114 106567
rect -55207 104041 -55190 104058
rect -55059 106553 -55042 106570
rect -54938 106544 -54921 106561
rect -55131 104027 -55114 104044
rect -55059 104030 -55042 104047
rect -53429 108900 -53367 108964
rect -53429 108400 -53367 108464
rect -53429 107900 -53367 107964
rect -53429 107400 -53367 107464
rect -53429 106900 -53367 106964
rect -53429 106400 -53367 106464
rect -53429 105900 -53367 105964
rect -53429 105400 -53367 105464
rect -54601 105107 -54557 105155
rect -54600 105020 -54556 105068
rect -54381 105106 -54337 105154
rect -54390 105004 -54344 105050
rect -54169 105107 -54125 105155
rect -54170 105013 -54126 105061
rect -53956 105103 -53902 105161
rect -53953 105015 -53907 105062
rect -53429 104900 -53367 104964
rect -54403 104592 -54340 104641
rect -54944 104015 -54919 104037
rect -54403 104392 -54340 104456
rect -54403 104192 -54340 104256
rect -54403 103992 -54340 104056
rect -54753 103726 -54705 103772
rect -54753 103526 -54705 103572
rect -54753 103326 -54705 103372
rect -54753 103126 -54705 103172
rect -54753 102926 -54705 102972
rect -54540 103729 -54492 103775
rect -54540 103529 -54492 103575
rect -54540 103329 -54492 103375
rect -54540 103129 -54492 103175
rect -54540 102929 -54492 102975
rect -54403 103792 -54340 103856
rect -54403 103592 -54340 103656
rect -54403 103392 -54340 103456
rect -54403 103192 -54340 103256
rect -54403 102992 -54340 103056
rect -54403 102792 -54340 102856
rect -54190 104592 -54127 104656
rect -54190 104392 -54127 104456
rect -54190 104192 -54127 104256
rect -54190 103992 -54127 104056
rect -54190 103792 -54127 103856
rect -54190 103592 -54127 103656
rect -54190 103392 -54127 103456
rect -54190 103192 -54127 103256
rect -54190 102992 -54127 103056
rect -54190 102792 -54127 102856
rect -53429 104400 -53367 104464
rect -53429 103900 -53367 103964
rect -53429 103400 -53367 103464
rect -53429 102900 -53367 102964
rect -53221 108900 -53159 108964
rect -53221 108400 -53159 108464
rect -53221 107900 -53159 107964
rect -53221 107400 -53159 107464
rect -53221 106900 -53159 106964
rect -53221 106400 -53159 106464
rect -53221 105900 -53159 105964
rect -53221 105400 -53159 105464
rect -53221 104900 -53159 104964
rect -53221 104400 -53159 104464
rect -53221 103900 -53159 103964
rect -53221 103400 -53159 103464
rect -53221 102900 -53159 102964
<< pdiffc >>
rect -53819 111334 -53751 111407
rect -53819 110834 -53751 110907
rect -53819 110334 -53751 110407
rect -53819 109834 -53751 109907
rect -53819 109334 -53751 109407
rect -53819 108834 -53751 108907
rect -53819 108334 -53751 108407
rect -53819 107834 -53751 107907
rect -53819 107334 -53751 107407
rect -53819 106834 -53751 106907
rect -53819 106334 -53751 106407
rect -54602 106135 -54535 106207
rect -54602 105935 -54535 106007
rect -54602 105735 -54535 105807
rect -54602 105535 -54535 105607
rect -54602 105335 -54535 105407
rect -54390 106134 -54322 106207
rect -54390 105934 -54322 106007
rect -54390 105734 -54322 105807
rect -54390 105534 -54322 105607
rect -54390 105334 -54322 105407
rect -54176 106134 -54108 106207
rect -54176 105934 -54108 106007
rect -54176 105734 -54108 105807
rect -54176 105534 -54108 105607
rect -54176 105334 -54108 105407
rect -53968 106134 -53900 106207
rect -53968 105934 -53900 106007
rect -53968 105734 -53900 105807
rect -53968 105534 -53900 105607
rect -53968 105334 -53900 105407
rect -53819 105834 -53751 105907
rect -53819 105334 -53751 105407
rect -53613 111334 -53545 111407
rect -53613 110834 -53545 110907
rect -53613 110334 -53545 110407
rect -53613 109834 -53545 109907
rect -53613 109334 -53545 109407
rect -53613 108834 -53545 108907
rect -53613 108334 -53545 108407
rect -53613 107834 -53545 107907
rect -53613 107334 -53545 107407
rect -53613 106834 -53545 106907
rect -53613 106334 -53545 106407
rect -53613 105834 -53545 105907
rect -53613 105334 -53545 105407
<< psubdiff >>
rect -55329 106559 -55253 106590
rect -55329 106509 -55317 106559
rect -55268 106509 -55253 106559
rect -55329 103782 -55253 106509
rect -53018 109133 -52940 109153
rect -55329 103750 -55251 103782
rect -55329 103692 -55322 103750
rect -55259 103692 -55251 103750
rect -55329 103664 -55251 103692
rect -55328 102640 -55251 103664
rect -53018 109093 -53005 109133
rect -52954 109093 -52940 109133
rect -53018 108633 -52940 109093
rect -53018 108593 -53005 108633
rect -52954 108593 -52940 108633
rect -53018 108133 -52940 108593
rect -53018 108093 -53005 108133
rect -52954 108093 -52940 108133
rect -53018 107633 -52940 108093
rect -53018 107593 -53005 107633
rect -52954 107593 -52940 107633
rect -53018 107133 -52940 107593
rect -53018 107093 -53005 107133
rect -52954 107093 -52940 107133
rect -53018 106633 -52940 107093
rect -53018 106593 -53005 106633
rect -52954 106593 -52940 106633
rect -53018 106133 -52940 106593
rect -53018 106093 -53005 106133
rect -52954 106093 -52940 106133
rect -53018 105633 -52940 106093
rect -53018 105593 -53005 105633
rect -52954 105593 -52940 105633
rect -53018 105133 -52940 105593
rect -53018 105093 -53005 105133
rect -52954 105093 -52940 105133
rect -53018 104633 -52940 105093
rect -53018 104593 -53005 104633
rect -52954 104593 -52940 104633
rect -53018 104133 -52940 104593
rect -53018 104093 -53005 104133
rect -52954 104093 -52940 104133
rect -53018 103633 -52940 104093
rect -53018 103593 -53005 103633
rect -52954 103593 -52940 103633
rect -53018 103133 -52940 103593
rect -53018 103093 -53005 103133
rect -52954 103093 -52940 103133
rect -53018 102640 -52940 103093
rect -55328 102633 -52940 102640
rect -55328 102631 -53005 102633
rect -55328 102592 -55313 102631
rect -55264 102627 -53005 102631
rect -55264 102592 -55009 102627
rect -55328 102588 -55009 102592
rect -54960 102625 -53005 102627
rect -54960 102588 -54687 102625
rect -55328 102585 -54687 102588
rect -54638 102585 -54187 102625
rect -54138 102585 -53687 102625
rect -53638 102585 -53187 102625
rect -53138 102593 -53005 102625
rect -52954 102593 -52940 102633
rect -53138 102585 -52940 102593
rect -55328 102576 -52940 102585
<< nsubdiff >>
rect -53955 111680 -53888 111681
rect -53957 111668 -53523 111680
rect -53957 111621 -53948 111668
rect -53901 111665 -53523 111668
rect -53901 111623 -53586 111665
rect -53538 111623 -53523 111665
rect -53901 111621 -53523 111623
rect -53957 111615 -53523 111621
rect -53955 111235 -53888 111615
rect -53955 111194 -53939 111235
rect -53902 111194 -53888 111235
rect -53955 110735 -53888 111194
rect -53955 110694 -53939 110735
rect -53902 110694 -53888 110735
rect -53955 110627 -53888 110694
rect -53955 110235 -53887 110627
rect -53955 110194 -53939 110235
rect -53902 110194 -53887 110235
rect -53955 110034 -53887 110194
rect -53954 109735 -53887 110034
rect -53954 109694 -53939 109735
rect -53902 109694 -53887 109735
rect -53954 109349 -53887 109694
rect -53954 109235 -53890 109349
rect -53954 109194 -53939 109235
rect -53902 109194 -53890 109235
rect -53954 108735 -53890 109194
rect -53954 108694 -53939 108735
rect -53902 108694 -53890 108735
rect -53954 108235 -53890 108694
rect -53954 108194 -53939 108235
rect -53902 108194 -53890 108235
rect -53954 107735 -53890 108194
rect -53954 107694 -53939 107735
rect -53902 107694 -53890 107735
rect -53954 107235 -53890 107694
rect -53954 107194 -53939 107235
rect -53902 107194 -53890 107235
rect -53954 106735 -53890 107194
rect -53954 106694 -53939 106735
rect -53902 106694 -53890 106735
rect -53954 106554 -53890 106694
rect -53953 106486 -53890 106554
rect -53953 106453 -53942 106486
rect -53909 106453 -53890 106486
rect -53953 106441 -53890 106453
rect -54580 106431 -53890 106441
rect -54580 106430 -54376 106431
rect -54580 106397 -54562 106430
rect -54529 106398 -54376 106430
rect -54343 106398 -54191 106431
rect -54158 106398 -54032 106431
rect -53999 106398 -53890 106431
rect -54529 106397 -53890 106398
rect -54580 106386 -53890 106397
<< psubdiffcont >>
rect -55317 106509 -55268 106559
rect -55322 103692 -55259 103750
rect -53005 109093 -52954 109133
rect -53005 108593 -52954 108633
rect -53005 108093 -52954 108133
rect -53005 107593 -52954 107633
rect -53005 107093 -52954 107133
rect -53005 106593 -52954 106633
rect -53005 106093 -52954 106133
rect -53005 105593 -52954 105633
rect -53005 105093 -52954 105133
rect -53005 104593 -52954 104633
rect -53005 104093 -52954 104133
rect -53005 103593 -52954 103633
rect -53005 103093 -52954 103133
rect -55313 102592 -55264 102631
rect -55009 102588 -54960 102627
rect -54687 102585 -54638 102625
rect -54187 102585 -54138 102625
rect -53687 102585 -53638 102625
rect -53187 102585 -53138 102625
rect -53005 102593 -52954 102633
<< nsubdiffcont >>
rect -53948 111621 -53901 111668
rect -53586 111623 -53538 111665
rect -53939 111194 -53902 111235
rect -53939 110694 -53902 110735
rect -53939 110194 -53902 110235
rect -53939 109694 -53902 109735
rect -53939 109194 -53902 109235
rect -53939 108694 -53902 108735
rect -53939 108194 -53902 108235
rect -53939 107694 -53902 107735
rect -53939 107194 -53902 107235
rect -53939 106694 -53902 106735
rect -53942 106453 -53909 106486
rect -54562 106397 -54529 106430
rect -54376 106398 -54343 106431
rect -54191 106398 -54158 106431
rect -54032 106398 -53999 106431
<< poly >>
rect -53733 111578 -53633 111601
rect -54518 106336 -54418 106349
rect -54518 106330 -54480 106336
rect -54520 106316 -54480 106330
rect -54453 106330 -54418 106336
rect -54453 106316 -53988 106330
rect -54520 106301 -53988 106316
rect -54518 106292 -54418 106301
rect -54089 106292 -53989 106301
rect -54518 105245 -54418 105291
rect -54089 105245 -53989 105291
rect -53346 109125 -53246 109148
rect -53733 105265 -53633 105289
rect -53733 105242 -53708 105265
rect -53648 105242 -53633 105265
rect -53733 105230 -53633 105242
rect -54518 105176 -54418 105210
rect -54088 105174 -53988 105208
rect -54518 104972 -54418 104997
rect -54088 104987 -53988 104995
rect -54518 104926 -54492 104972
rect -54445 104926 -54418 104972
rect -54518 104906 -54418 104926
rect -54089 104933 -53988 104987
rect -54089 104898 -54060 104933
rect -54020 104898 -53988 104933
rect -54089 104875 -53988 104898
rect -54317 104755 -54217 104780
rect -54678 103941 -54578 103949
rect -54678 103913 -54656 103941
rect -54597 103913 -54578 103941
rect -54678 103894 -54578 103913
rect -54678 102715 -54578 102893
rect -54317 102715 -54217 102753
rect -53346 102715 -53246 102836
rect -54678 102679 -53246 102715
<< polycont >>
rect -54480 106316 -54453 106336
rect -53708 105242 -53648 105265
rect -54492 104926 -54445 104972
rect -54060 104898 -54020 104933
rect -54656 103913 -54597 103941
<< ndiffres >>
rect -55217 106588 -55180 106590
rect -55217 106557 -55212 106588
rect -55185 106557 -55180 106588
rect -55217 104421 -55180 106557
rect -55141 106574 -55104 106591
rect -55141 106543 -55136 106574
rect -55109 106543 -55104 106574
rect -55217 104065 -55181 104421
rect -55217 104034 -55212 104065
rect -55185 104034 -55181 104065
rect -55217 104028 -55181 104034
rect -55141 104407 -55104 106543
rect -55069 106577 -55032 106594
rect -55069 106546 -55064 106577
rect -55037 106546 -55032 106577
rect -55069 104410 -55032 106546
rect -54948 106568 -54911 106572
rect -54948 106537 -54943 106568
rect -54916 106537 -54911 106568
rect -55141 104051 -55105 104407
rect -55141 104020 -55136 104051
rect -55109 104020 -55105 104051
rect -55141 104014 -55105 104020
rect -55069 104054 -55033 104410
rect -55069 104023 -55064 104054
rect -55037 104023 -55033 104054
rect -55069 104017 -55033 104023
rect -54948 104401 -54911 106537
rect -54948 104043 -54912 104401
rect -54948 104012 -54944 104043
rect -54917 104037 -54912 104043
rect -54919 104015 -54912 104037
rect -54917 104012 -54912 104015
rect -54948 104006 -54912 104012
<< locali >>
rect -66599 125061 -65639 125392
rect -66599 124993 -51996 125061
rect -66599 124302 -66428 124993
rect -65899 124302 -51996 124993
rect -66599 124155 -51996 124302
rect -66599 123870 -65639 124155
rect -59529 115127 -53654 115302
rect -59529 114718 -59190 115127
rect -58652 114718 -53654 115127
rect -59529 114528 -53654 114718
rect -59079 114527 -59057 114528
rect -53704 112119 -53654 114528
rect -53850 111989 -53654 112119
rect -53850 111891 -53655 111989
rect -53955 111680 -53888 111681
rect -53847 111680 -53797 111891
rect -53957 111668 -53523 111680
rect -53957 111621 -53948 111668
rect -53901 111665 -53523 111668
rect -53901 111623 -53586 111665
rect -53538 111623 -53523 111665
rect -53901 111621 -53523 111623
rect -53957 111615 -53523 111621
rect -53955 111235 -53888 111615
rect -53807 111418 -53762 111615
rect -53828 111407 -53741 111418
rect -53828 111334 -53819 111407
rect -53751 111334 -53741 111407
rect -53828 111326 -53741 111334
rect -53622 111407 -53535 111417
rect -53622 111334 -53613 111407
rect -53545 111334 -53535 111407
rect -53622 111325 -53535 111334
rect -53955 111194 -53939 111235
rect -53902 111194 -53888 111235
rect -53955 110735 -53888 111194
rect -53828 110907 -53741 110918
rect -53828 110834 -53819 110907
rect -53751 110834 -53741 110907
rect -53828 110826 -53741 110834
rect -53622 110907 -53535 110917
rect -53622 110834 -53613 110907
rect -53545 110834 -53535 110907
rect -53622 110825 -53535 110834
rect -53955 110694 -53939 110735
rect -53902 110694 -53888 110735
rect -53955 110627 -53888 110694
rect -53955 110235 -53887 110627
rect -53828 110407 -53741 110418
rect -53828 110334 -53819 110407
rect -53751 110334 -53741 110407
rect -53828 110326 -53741 110334
rect -53622 110407 -53535 110417
rect -53622 110334 -53613 110407
rect -53545 110334 -53535 110407
rect -53622 110325 -53535 110334
rect -53955 110194 -53939 110235
rect -53902 110194 -53887 110235
rect -53955 110034 -53887 110194
rect -53954 109735 -53887 110034
rect -53828 109907 -53741 109918
rect -53828 109834 -53819 109907
rect -53751 109834 -53741 109907
rect -53828 109826 -53741 109834
rect -53622 109907 -53535 109917
rect -53622 109834 -53613 109907
rect -53545 109834 -53535 109907
rect -53622 109825 -53535 109834
rect -53954 109694 -53939 109735
rect -53902 109694 -53887 109735
rect -53954 109349 -53887 109694
rect -53828 109407 -53741 109418
rect -53954 109235 -53890 109349
rect -53828 109334 -53819 109407
rect -53751 109334 -53741 109407
rect -53828 109326 -53741 109334
rect -53622 109413 -53535 109417
rect -53059 109413 -51996 124155
rect -53622 109407 -51996 109413
rect -53622 109334 -53613 109407
rect -53545 109334 -51996 109407
rect -53622 109329 -51996 109334
rect -53622 109325 -53535 109329
rect -53954 109194 -53939 109235
rect -53902 109194 -53890 109235
rect -53954 108735 -53890 109194
rect -53418 108978 -53378 109329
rect -53018 109133 -52940 109153
rect -53018 109093 -53005 109133
rect -52954 109093 -52940 109133
rect -53441 108964 -53354 108978
rect -53828 108907 -53741 108918
rect -53828 108834 -53819 108907
rect -53751 108834 -53741 108907
rect -53828 108826 -53741 108834
rect -53622 108907 -53535 108917
rect -53622 108834 -53613 108907
rect -53545 108834 -53535 108907
rect -53441 108900 -53429 108964
rect -53367 108900 -53354 108964
rect -53441 108886 -53354 108900
rect -53233 108964 -53146 108978
rect -53233 108900 -53221 108964
rect -53159 108900 -53146 108964
rect -53233 108886 -53146 108900
rect -53622 108825 -53535 108834
rect -53954 108694 -53939 108735
rect -53902 108694 -53890 108735
rect -53954 108235 -53890 108694
rect -53018 108633 -52940 109093
rect -53018 108593 -53005 108633
rect -52954 108593 -52940 108633
rect -53441 108464 -53354 108478
rect -53828 108407 -53741 108418
rect -53828 108334 -53819 108407
rect -53751 108334 -53741 108407
rect -53828 108326 -53741 108334
rect -53622 108407 -53535 108417
rect -53622 108334 -53613 108407
rect -53545 108334 -53535 108407
rect -53441 108400 -53429 108464
rect -53367 108400 -53354 108464
rect -53441 108386 -53354 108400
rect -53233 108464 -53146 108478
rect -53233 108400 -53221 108464
rect -53159 108400 -53146 108464
rect -53233 108386 -53146 108400
rect -53622 108325 -53535 108334
rect -53954 108194 -53939 108235
rect -53902 108194 -53890 108235
rect -53954 107735 -53890 108194
rect -53018 108133 -52940 108593
rect -53018 108093 -53005 108133
rect -52954 108093 -52940 108133
rect -53441 107964 -53354 107978
rect -53828 107907 -53741 107918
rect -53828 107834 -53819 107907
rect -53751 107834 -53741 107907
rect -53828 107826 -53741 107834
rect -53622 107907 -53535 107917
rect -53622 107834 -53613 107907
rect -53545 107834 -53535 107907
rect -53441 107900 -53429 107964
rect -53367 107900 -53354 107964
rect -53441 107886 -53354 107900
rect -53233 107964 -53146 107978
rect -53233 107900 -53221 107964
rect -53159 107900 -53146 107964
rect -53233 107886 -53146 107900
rect -53622 107825 -53535 107834
rect -53954 107694 -53939 107735
rect -53902 107694 -53890 107735
rect -61604 107096 -55561 107501
rect -53954 107235 -53890 107694
rect -53018 107633 -52940 108093
rect -53018 107593 -53005 107633
rect -52954 107593 -52940 107633
rect -53441 107464 -53354 107478
rect -53828 107407 -53741 107418
rect -53828 107334 -53819 107407
rect -53751 107334 -53741 107407
rect -53828 107326 -53741 107334
rect -53622 107407 -53535 107417
rect -53622 107334 -53613 107407
rect -53545 107334 -53535 107407
rect -53441 107400 -53429 107464
rect -53367 107400 -53354 107464
rect -53441 107386 -53354 107400
rect -53233 107464 -53146 107478
rect -53233 107400 -53221 107464
rect -53159 107400 -53146 107464
rect -53233 107386 -53146 107400
rect -53622 107325 -53535 107334
rect -53954 107194 -53939 107235
rect -53902 107194 -53890 107235
rect -61604 106974 -54680 107096
rect -61604 106958 -55561 106974
rect -61559 53027 -61219 106958
rect -54734 106876 -54680 106974
rect -55527 106816 -54790 106819
rect -55631 106810 -54790 106816
rect -55631 106781 -54828 106810
rect -54794 106781 -54790 106810
rect -55631 106757 -54790 106781
rect -55631 106728 -54830 106757
rect -54796 106728 -54790 106757
rect -55631 106719 -54790 106728
rect -54733 106761 -54684 106876
rect -54733 106729 -54723 106761
rect -54692 106729 -54684 106761
rect -54733 106719 -54684 106729
rect -53954 106735 -53890 107194
rect -53018 107133 -52940 107593
rect -53018 107093 -53005 107133
rect -52954 107093 -52940 107133
rect -53441 106964 -53354 106978
rect -53828 106907 -53741 106918
rect -53828 106834 -53819 106907
rect -53751 106834 -53741 106907
rect -53828 106826 -53741 106834
rect -53622 106907 -53535 106917
rect -53622 106834 -53613 106907
rect -53545 106834 -53535 106907
rect -53441 106900 -53429 106964
rect -53367 106900 -53354 106964
rect -53441 106886 -53354 106900
rect -53233 106964 -53146 106978
rect -53233 106900 -53221 106964
rect -53159 106900 -53146 106964
rect -53233 106886 -53146 106900
rect -53622 106825 -53535 106834
rect -56606 106594 -56229 106603
rect -55631 106594 -55452 106719
rect -53954 106694 -53939 106735
rect -53902 106694 -53890 106735
rect -55210 106630 -54539 106656
rect -56609 106443 -55449 106594
rect -55210 106590 -55188 106630
rect -55067 106594 -55033 106596
rect -55139 106591 -55105 106592
rect -55329 106559 -55253 106590
rect -55329 106509 -55317 106559
rect -55268 106509 -55253 106559
rect -55215 106581 -55180 106590
rect -55215 106564 -55207 106581
rect -55190 106564 -55180 106581
rect -55215 106554 -55180 106564
rect -55214 106546 -55180 106554
rect -55139 106583 -55104 106591
rect -55067 106583 -55032 106594
rect -55139 106570 -55032 106583
rect -55139 106567 -55059 106570
rect -55139 106550 -55131 106567
rect -55114 106553 -55059 106567
rect -55042 106553 -55032 106570
rect -54948 106565 -54911 106572
rect -55114 106550 -55032 106553
rect -55139 106548 -55032 106550
rect -55139 106540 -55104 106548
rect -55067 106543 -55032 106548
rect -55138 106532 -55104 106540
rect -55066 106535 -55032 106543
rect -55000 106561 -54911 106565
rect -55000 106544 -54938 106561
rect -54921 106544 -54911 106561
rect -55000 106543 -54911 106544
rect -62501 52846 -61219 53027
rect -62501 52494 -62103 52846
rect -61490 52494 -61219 52846
rect -62501 52420 -61219 52494
rect -62501 52380 -61241 52420
rect -56606 31242 -56229 106443
rect -55329 103782 -55253 106509
rect -55218 104058 -55172 104079
rect -55218 104041 -55207 104058
rect -55190 104047 -55172 104058
rect -55150 104047 -55096 104065
rect -55190 104044 -55096 104047
rect -55190 104041 -55131 104044
rect -55218 104027 -55131 104041
rect -55114 104027 -55096 104044
rect -55147 104008 -55096 104027
rect -55078 104047 -55024 104068
rect -55078 104030 -55059 104047
rect -55042 104030 -55024 104047
rect -55078 104019 -55024 104030
rect -55075 104007 -55024 104019
rect -55000 104007 -54975 106543
rect -54949 106535 -54911 106543
rect -54570 106441 -54539 106630
rect -53954 106554 -53890 106694
rect -53953 106486 -53890 106554
rect -53953 106453 -53942 106486
rect -53909 106453 -53890 106486
rect -53018 106633 -52940 107093
rect -53018 106593 -53005 106633
rect -52954 106593 -52940 106633
rect -53953 106441 -53890 106453
rect -54580 106431 -53890 106441
rect -54580 106430 -54376 106431
rect -54580 106397 -54562 106430
rect -54529 106398 -54376 106430
rect -54343 106398 -54191 106431
rect -54158 106398 -54032 106431
rect -53999 106398 -53890 106431
rect -53441 106464 -53354 106478
rect -54529 106397 -53890 106398
rect -54580 106386 -53890 106397
rect -53828 106407 -53741 106418
rect -54518 106336 -54418 106343
rect -54518 106330 -54480 106336
rect -54602 106316 -54480 106330
rect -54453 106316 -54418 106336
rect -54602 106300 -54418 106316
rect -54602 106218 -54540 106300
rect -54518 106299 -54418 106300
rect -54386 106218 -54327 106386
rect -54171 106218 -54113 106386
rect -53828 106334 -53819 106407
rect -53751 106334 -53741 106407
rect -53828 106326 -53741 106334
rect -53622 106407 -53535 106417
rect -53622 106334 -53613 106407
rect -53545 106334 -53535 106407
rect -53441 106400 -53429 106464
rect -53367 106400 -53354 106464
rect -53441 106386 -53354 106400
rect -53233 106464 -53146 106478
rect -53233 106400 -53221 106464
rect -53159 106400 -53146 106464
rect -53233 106386 -53146 106400
rect -53622 106325 -53535 106334
rect -54611 106207 -54524 106218
rect -54611 106135 -54602 106207
rect -54535 106135 -54524 106207
rect -54611 106126 -54524 106135
rect -54400 106207 -54313 106218
rect -54400 106134 -54390 106207
rect -54322 106134 -54313 106207
rect -54400 106126 -54313 106134
rect -54185 106207 -54098 106218
rect -54185 106134 -54176 106207
rect -54108 106134 -54098 106207
rect -54185 106126 -54098 106134
rect -53978 106207 -53891 106218
rect -53978 106134 -53968 106207
rect -53900 106134 -53891 106207
rect -53978 106126 -53891 106134
rect -53018 106133 -52940 106593
rect -53018 106093 -53005 106133
rect -52954 106093 -52940 106133
rect -54611 106007 -54524 106018
rect -54611 105935 -54602 106007
rect -54535 105935 -54524 106007
rect -54611 105926 -54524 105935
rect -54400 106007 -54313 106018
rect -54400 105934 -54390 106007
rect -54322 105934 -54313 106007
rect -54400 105926 -54313 105934
rect -54185 106007 -54098 106018
rect -54185 105934 -54176 106007
rect -54108 105934 -54098 106007
rect -54185 105926 -54098 105934
rect -53978 106007 -53891 106018
rect -53978 105934 -53968 106007
rect -53900 105934 -53891 106007
rect -53978 105926 -53891 105934
rect -53441 105964 -53354 105978
rect -53828 105907 -53741 105918
rect -53828 105834 -53819 105907
rect -53751 105834 -53741 105907
rect -53828 105826 -53741 105834
rect -53622 105907 -53535 105917
rect -53622 105834 -53613 105907
rect -53545 105834 -53535 105907
rect -53441 105900 -53429 105964
rect -53367 105900 -53354 105964
rect -53441 105886 -53354 105900
rect -53233 105964 -53146 105978
rect -53233 105900 -53221 105964
rect -53159 105900 -53146 105964
rect -53233 105886 -53146 105900
rect -53622 105825 -53535 105834
rect -54611 105807 -54524 105818
rect -54611 105735 -54602 105807
rect -54535 105735 -54524 105807
rect -54611 105726 -54524 105735
rect -54400 105807 -54313 105818
rect -54400 105734 -54390 105807
rect -54322 105734 -54313 105807
rect -54400 105726 -54313 105734
rect -54185 105807 -54098 105818
rect -54185 105734 -54176 105807
rect -54108 105734 -54098 105807
rect -54185 105726 -54098 105734
rect -53978 105807 -53891 105818
rect -53978 105734 -53968 105807
rect -53900 105734 -53891 105807
rect -53978 105726 -53891 105734
rect -53018 105633 -52940 106093
rect -54611 105607 -54524 105618
rect -54611 105535 -54602 105607
rect -54535 105535 -54524 105607
rect -54611 105526 -54524 105535
rect -54400 105607 -54313 105618
rect -54400 105534 -54390 105607
rect -54322 105534 -54313 105607
rect -54400 105526 -54313 105534
rect -54185 105607 -54098 105618
rect -54185 105534 -54176 105607
rect -54108 105534 -54098 105607
rect -54185 105526 -54098 105534
rect -53978 105607 -53891 105618
rect -53978 105534 -53968 105607
rect -53900 105534 -53891 105607
rect -53978 105526 -53891 105534
rect -53018 105593 -53005 105633
rect -52954 105593 -52940 105633
rect -53441 105464 -53354 105478
rect -54611 105407 -54524 105418
rect -54611 105335 -54602 105407
rect -54535 105335 -54524 105407
rect -54611 105326 -54524 105335
rect -54400 105407 -54313 105418
rect -54400 105334 -54390 105407
rect -54322 105334 -54313 105407
rect -54400 105326 -54313 105334
rect -54186 105407 -54099 105418
rect -54186 105334 -54176 105407
rect -54108 105334 -54099 105407
rect -54186 105326 -54099 105334
rect -53978 105407 -53891 105418
rect -53978 105334 -53968 105407
rect -53900 105334 -53891 105407
rect -53978 105326 -53891 105334
rect -53828 105407 -53741 105418
rect -53828 105334 -53819 105407
rect -53751 105334 -53741 105407
rect -53828 105326 -53741 105334
rect -53622 105407 -53535 105417
rect -53622 105334 -53613 105407
rect -53545 105334 -53535 105407
rect -53441 105400 -53429 105464
rect -53367 105400 -53354 105464
rect -53441 105386 -53354 105400
rect -53233 105464 -53146 105478
rect -53233 105400 -53221 105464
rect -53159 105400 -53146 105464
rect -53233 105386 -53146 105400
rect -54601 105165 -54555 105326
rect -53964 105275 -53897 105326
rect -53622 105325 -53535 105334
rect -53733 105275 -53633 105284
rect -53964 105265 -53633 105275
rect -53964 105242 -53708 105265
rect -53648 105242 -53633 105265
rect -53964 105241 -53633 105242
rect -54613 105155 -54547 105165
rect -54613 105107 -54601 105155
rect -54557 105107 -54547 105155
rect -54613 105094 -54547 105107
rect -54393 105154 -54327 105165
rect -54393 105106 -54381 105154
rect -54337 105106 -54327 105154
rect -54393 105095 -54327 105106
rect -54183 105155 -54117 105163
rect -54183 105107 -54169 105155
rect -54125 105107 -54117 105155
rect -53964 105161 -53897 105241
rect -53733 105230 -53633 105241
rect -53964 105125 -53956 105161
rect -54183 105092 -54117 105107
rect -53963 105103 -53956 105125
rect -53902 105103 -53897 105161
rect -53963 105092 -53897 105103
rect -53018 105133 -52940 105593
rect -53018 105093 -53005 105133
rect -52954 105093 -52940 105133
rect -54613 105068 -54547 105076
rect -54613 105020 -54600 105068
rect -54556 105020 -54547 105068
rect -54613 105005 -54547 105020
rect -54405 105061 -54329 105065
rect -54183 105061 -54117 105074
rect -54405 105050 -54170 105061
rect -54405 105004 -54390 105050
rect -54344 105013 -54170 105050
rect -54126 105013 -54117 105061
rect -54344 105004 -54117 105013
rect -53963 105062 -53897 105075
rect -53963 105015 -53953 105062
rect -53907 105015 -53897 105062
rect -53963 105004 -53897 105015
rect -54405 105003 -54117 105004
rect -54405 105001 -54123 105003
rect -54511 104972 -54426 104986
rect -54511 104926 -54492 104972
rect -54445 104926 -54426 104972
rect -54511 104907 -54426 104926
rect -54405 104755 -54329 105001
rect -53441 104964 -53354 104978
rect -54070 104933 -54010 104955
rect -54070 104898 -54060 104933
rect -54020 104898 -54010 104933
rect -54070 104852 -54010 104898
rect -53441 104900 -53429 104964
rect -53367 104900 -53354 104964
rect -53441 104886 -53354 104900
rect -53233 104964 -53146 104978
rect -53233 104900 -53221 104964
rect -53159 104900 -53146 104964
rect -53233 104886 -53146 104900
rect -54070 104820 -54058 104852
rect -54020 104820 -54010 104852
rect -54070 104812 -54010 104820
rect -54412 104641 -54330 104755
rect -54412 104592 -54403 104641
rect -54340 104592 -54330 104641
rect -54412 104583 -54330 104592
rect -54201 104656 -54119 104668
rect -54201 104592 -54190 104656
rect -54127 104592 -54119 104656
rect -54201 104583 -54119 104592
rect -53018 104633 -52940 105093
rect -53018 104593 -53005 104633
rect -52954 104593 -52940 104633
rect -54412 104456 -54330 104468
rect -54412 104392 -54403 104456
rect -54340 104392 -54330 104456
rect -54412 104383 -54330 104392
rect -54201 104456 -54119 104468
rect -54201 104392 -54190 104456
rect -54127 104392 -54119 104456
rect -54201 104383 -54119 104392
rect -53441 104464 -53354 104478
rect -53441 104400 -53429 104464
rect -53367 104400 -53354 104464
rect -53441 104386 -53354 104400
rect -53233 104464 -53146 104478
rect -53233 104400 -53221 104464
rect -53159 104400 -53146 104464
rect -53233 104386 -53146 104400
rect -54412 104256 -54330 104268
rect -54412 104192 -54403 104256
rect -54340 104192 -54330 104256
rect -54412 104183 -54330 104192
rect -54201 104256 -54119 104268
rect -54201 104192 -54190 104256
rect -54127 104192 -54119 104256
rect -54201 104183 -54119 104192
rect -53018 104133 -52940 104593
rect -53018 104093 -53005 104133
rect -52954 104093 -52940 104133
rect -54412 104056 -54330 104068
rect -55075 103987 -54975 104007
rect -54955 104037 -54911 104042
rect -54955 104015 -54944 104037
rect -54919 104015 -54911 104037
rect -54955 104007 -54911 104015
rect -54955 103968 -54705 104007
rect -54412 103992 -54403 104056
rect -54340 103992 -54330 104056
rect -54412 103983 -54330 103992
rect -54201 104056 -54119 104068
rect -54201 103992 -54190 104056
rect -54127 103992 -54119 104056
rect -54201 103983 -54119 103992
rect -54743 103942 -54705 103968
rect -53441 103964 -53354 103978
rect -54678 103942 -54578 103945
rect -54743 103941 -54578 103942
rect -54743 103913 -54656 103941
rect -54597 103913 -54578 103941
rect -54743 103897 -54578 103913
rect -53441 103900 -53429 103964
rect -53367 103900 -53354 103964
rect -54743 103784 -54705 103897
rect -53441 103886 -53354 103900
rect -53233 103964 -53146 103978
rect -53233 103900 -53221 103964
rect -53159 103900 -53146 103964
rect -53233 103886 -53146 103900
rect -54412 103856 -54330 103868
rect -54412 103792 -54403 103856
rect -54340 103792 -54330 103856
rect -55329 103750 -55251 103782
rect -55329 103692 -55322 103750
rect -55259 103692 -55251 103750
rect -54766 103772 -54692 103784
rect -54766 103726 -54753 103772
rect -54705 103726 -54692 103772
rect -54766 103712 -54692 103726
rect -54553 103775 -54479 103788
rect -54412 103783 -54330 103792
rect -54201 103856 -54119 103868
rect -54201 103792 -54190 103856
rect -54127 103792 -54119 103856
rect -54201 103783 -54119 103792
rect -54553 103729 -54540 103775
rect -54492 103729 -54479 103775
rect -54553 103715 -54479 103729
rect -55329 103664 -55251 103692
rect -55328 102640 -55251 103664
rect -54412 103656 -54330 103668
rect -54412 103592 -54403 103656
rect -54340 103592 -54330 103656
rect -54766 103572 -54692 103585
rect -54766 103526 -54753 103572
rect -54705 103526 -54692 103572
rect -54766 103512 -54692 103526
rect -54553 103575 -54479 103588
rect -54412 103583 -54330 103592
rect -54201 103656 -54119 103668
rect -54201 103592 -54190 103656
rect -54127 103592 -54119 103656
rect -54201 103583 -54119 103592
rect -53018 103633 -52940 104093
rect -53018 103593 -53005 103633
rect -52954 103593 -52940 103633
rect -54553 103529 -54540 103575
rect -54492 103529 -54479 103575
rect -54553 103515 -54479 103529
rect -54412 103456 -54330 103468
rect -54412 103392 -54403 103456
rect -54340 103392 -54330 103456
rect -54766 103372 -54692 103385
rect -54766 103326 -54753 103372
rect -54705 103326 -54692 103372
rect -54766 103312 -54692 103326
rect -54553 103375 -54479 103388
rect -54412 103383 -54330 103392
rect -54201 103456 -54119 103468
rect -54201 103392 -54190 103456
rect -54127 103392 -54119 103456
rect -54201 103383 -54119 103392
rect -53441 103464 -53354 103478
rect -53441 103400 -53429 103464
rect -53367 103400 -53354 103464
rect -53441 103386 -53354 103400
rect -53233 103464 -53146 103478
rect -53233 103400 -53221 103464
rect -53159 103400 -53146 103464
rect -53233 103386 -53146 103400
rect -54553 103329 -54540 103375
rect -54492 103329 -54479 103375
rect -54553 103315 -54479 103329
rect -54412 103256 -54330 103268
rect -54412 103192 -54403 103256
rect -54340 103192 -54330 103256
rect -54766 103172 -54692 103185
rect -54766 103126 -54753 103172
rect -54705 103126 -54692 103172
rect -54766 103112 -54692 103126
rect -54553 103175 -54479 103188
rect -54412 103183 -54330 103192
rect -54201 103256 -54119 103268
rect -54201 103192 -54190 103256
rect -54127 103192 -54119 103256
rect -54201 103183 -54119 103192
rect -54553 103129 -54540 103175
rect -54492 103129 -54479 103175
rect -54553 103115 -54479 103129
rect -53018 103133 -52940 103593
rect -53018 103093 -53005 103133
rect -52954 103093 -52940 103133
rect -54412 103056 -54330 103068
rect -54412 102992 -54403 103056
rect -54340 102992 -54330 103056
rect -54768 102972 -54693 102984
rect -54768 102926 -54753 102972
rect -54705 102926 -54693 102972
rect -54768 102910 -54693 102926
rect -54555 102975 -54480 102987
rect -54412 102983 -54330 102992
rect -54201 103056 -54119 103068
rect -54201 102992 -54190 103056
rect -54127 102992 -54119 103056
rect -54201 102983 -54119 102992
rect -54555 102929 -54540 102975
rect -54492 102929 -54480 102975
rect -54555 102913 -54480 102929
rect -53441 102964 -53354 102978
rect -54546 102640 -54484 102913
rect -53441 102900 -53429 102964
rect -53367 102900 -53354 102964
rect -53441 102886 -53354 102900
rect -53233 102964 -53146 102978
rect -53233 102900 -53221 102964
rect -53159 102956 -53146 102964
rect -53018 102956 -52940 103093
rect -53159 102910 -52940 102956
rect -53159 102900 -53146 102910
rect -53233 102886 -53146 102900
rect -54412 102856 -54330 102868
rect -54412 102792 -54403 102856
rect -54340 102792 -54330 102856
rect -54412 102783 -54330 102792
rect -54201 102856 -54119 102868
rect -54201 102792 -54190 102856
rect -54127 102792 -54119 102856
rect -54201 102783 -54119 102792
rect -54190 102640 -54129 102783
rect -53018 102640 -52940 102910
rect -55328 102633 -52940 102640
rect -55328 102631 -53005 102633
rect -55328 102592 -55313 102631
rect -55264 102627 -53005 102631
rect -55264 102592 -55009 102627
rect -55328 102588 -55009 102592
rect -54960 102625 -53005 102627
rect -54960 102588 -54687 102625
rect -55328 102585 -54687 102588
rect -54638 102585 -54187 102625
rect -54138 102585 -53687 102625
rect -53638 102585 -53187 102625
rect -53138 102593 -53005 102625
rect -52954 102593 -52940 102633
rect -53138 102585 -52940 102593
rect -55328 102576 -52940 102585
rect -53717 102322 -53613 102576
rect -53859 78813 -53132 102322
rect -54171 78790 -52613 78813
rect -54179 78513 -52613 78790
rect -54179 77730 -53818 78513
rect -52874 77730 -52613 78513
rect -54179 77469 -52613 77730
rect -54171 77454 -52613 77469
rect -57328 31116 -56157 31242
rect -57328 30863 -56998 31116
rect -56361 30863 -56157 31116
rect -57328 30779 -56157 30863
<< viali >>
rect -66428 124302 -65899 124993
rect -62308 114712 -61770 115121
rect -61357 114707 -60819 115116
rect -60545 114714 -60007 115123
rect -59190 114718 -58652 115127
rect -54828 106781 -54794 106810
rect -54830 106728 -54796 106757
rect -54723 106729 -54692 106761
rect -62103 52494 -61490 52846
rect -54482 104935 -54459 104961
rect -54058 104820 -54020 104852
rect -53818 77730 -52874 78513
rect -56998 30863 -56361 31116
<< metal1 >>
rect -66599 124993 -65639 125392
rect -66599 124302 -66428 124993
rect -65899 124302 -65639 124993
rect -66599 123870 -65639 124302
rect -62752 115127 -58419 115300
rect -62752 115123 -59190 115127
rect -62752 115121 -60545 115123
rect -62752 114712 -62308 115121
rect -61770 115116 -60545 115121
rect -61770 114712 -61357 115116
rect -62752 114707 -61357 114712
rect -60819 114712 -60545 115116
rect -60007 114718 -59190 115123
rect -58652 114718 -58419 115127
rect -60007 114712 -58419 114718
rect -60819 114707 -58419 114712
rect -62752 114527 -58419 114707
rect -54839 106810 -54790 106819
rect -54839 106781 -54828 106810
rect -54794 106781 -54790 106810
rect -54839 106757 -54790 106781
rect -54839 106728 -54830 106757
rect -54796 106728 -54790 106757
rect -54839 104861 -54790 106728
rect -54733 106761 -54684 106771
rect -54733 106729 -54723 106761
rect -54692 106729 -54684 106761
rect -54733 104976 -54684 106729
rect -54733 104961 -54443 104976
rect -54733 104935 -54482 104961
rect -54459 104935 -54443 104961
rect -54733 104925 -54443 104935
rect -54839 104852 -54010 104861
rect -54839 104820 -54058 104852
rect -54020 104820 -54010 104852
rect -54839 104812 -54010 104820
rect -54179 78513 -52628 78790
rect -54179 77730 -53818 78513
rect -52874 77730 -52628 78513
rect -54179 77469 -52628 77730
rect -62482 52846 -61177 53038
rect -62482 52494 -62103 52846
rect -61490 52494 -61177 52846
rect -62482 52357 -61177 52494
rect -57328 31116 -56157 31242
rect -57328 30863 -56998 31116
rect -56361 30863 -56157 31116
rect -57328 30779 -56157 30863
<< via1 >>
rect -66428 124302 -65899 124993
rect -62308 114712 -61770 115121
rect -61357 114707 -60819 115116
rect -60545 114714 -60007 115121
rect -60545 114712 -60007 114714
rect -53818 77730 -52874 78513
rect -62103 52494 -61490 52846
rect -56998 30863 -56361 31116
<< metal2 >>
rect -66599 124993 -65639 125392
rect -66599 124302 -66428 124993
rect -65899 124302 -65639 124993
rect -66599 123870 -65639 124302
rect -62752 115121 -58419 115300
rect -62752 114712 -62308 115121
rect -61770 115116 -60545 115121
rect -61770 114712 -61357 115116
rect -62752 114707 -61357 114712
rect -60819 114712 -60545 115116
rect -60007 114712 -58419 115121
rect -60819 114707 -58419 114712
rect -62752 114527 -58419 114707
rect -54179 78513 -52628 78790
rect -54179 77730 -53818 78513
rect -52874 77730 -52628 78513
rect -54179 77469 -52628 77730
rect -62482 52846 -61177 53038
rect -62482 52494 -62103 52846
rect -61490 52494 -61177 52846
rect -62482 52357 -61177 52494
rect -57328 31116 -56157 31242
rect -57328 30863 -56998 31116
rect -56361 30863 -56157 31116
rect -57328 30779 -56157 30863
<< via2 >>
rect -66428 124302 -65899 124993
rect -62308 114712 -61770 115121
rect -61357 114707 -60819 115116
rect -60545 114712 -60007 115121
rect -53818 77730 -52874 78513
rect -62103 52494 -61490 52846
rect -56998 30863 -56361 31116
<< metal3 >>
rect -66681 136547 -66218 137753
rect -66681 135094 -66205 136547
rect -66610 125392 -66205 135094
rect -66610 124993 -65639 125392
rect -66610 124302 -66428 124993
rect -65899 124302 -65639 124993
rect -66610 123890 -65639 124302
rect -66599 123870 -65639 123890
rect -66595 115300 -64884 115309
rect -66595 115121 -58419 115300
rect -66595 114712 -62308 115121
rect -61770 115116 -60545 115121
rect -61770 114712 -61357 115116
rect -66595 114707 -61357 114712
rect -60819 114712 -60545 115116
rect -60007 114712 -58419 115121
rect -60819 114707 -58419 114712
rect -66595 114527 -58419 114707
rect -66595 114526 -64884 114527
rect -54171 78513 -52613 78813
rect -54171 78012 -53818 78513
rect -66729 77730 -53818 78012
rect -52874 77730 -52613 78513
rect -66729 77466 -52613 77730
rect -54171 77454 -52613 77466
rect -64339 52846 -61229 53038
rect -64339 52845 -62103 52846
rect -67009 52494 -62103 52845
rect -61490 52494 -61229 52846
rect -67009 52376 -61229 52494
rect -64339 52357 -61229 52376
rect -64716 31252 -61805 31254
rect -66924 31245 -61805 31252
rect -59455 31245 -56187 31248
rect -66924 31116 -56187 31245
rect -66924 30863 -56998 31116
rect -56361 30863 -56187 31116
rect -66924 30785 -56187 30863
rect -66924 30783 -64013 30785
rect -62229 30779 -56187 30785
rect -62229 30777 -56980 30779
rect -62229 30776 -59318 30777
<< labels >>
rlabel locali -53760 111645 -53760 111645 1 vdd
rlabel locali -53403 109371 -53403 109371 1 out
rlabel locali -53890 102601 -53890 102601 1 vss
rlabel locali -54044 104946 -54044 104946 1 in2
rlabel locali -54471 104979 -54471 104979 1 in1
<< end >>
